
module REG_ID ( clk, in, instr );
  input [31:0] in;
  output [31:0] instr;
  input clk;


  DFF_X1 instr_reg_31_ ( .D(in[31]), .CK(clk), .Q(instr[31]) );
  DFF_X1 instr_reg_30_ ( .D(in[30]), .CK(clk), .Q(instr[30]) );
  DFF_X1 instr_reg_29_ ( .D(in[29]), .CK(clk), .Q(instr[29]) );
  DFF_X1 instr_reg_28_ ( .D(in[28]), .CK(clk), .Q(instr[28]) );
  DFF_X1 instr_reg_27_ ( .D(in[27]), .CK(clk), .Q(instr[27]) );
  DFF_X1 instr_reg_26_ ( .D(in[26]), .CK(clk), .Q(instr[26]) );
  DFF_X1 instr_reg_25_ ( .D(in[25]), .CK(clk), .Q(instr[25]) );
  DFF_X1 instr_reg_24_ ( .D(in[24]), .CK(clk), .Q(instr[24]) );
  DFF_X1 instr_reg_23_ ( .D(in[23]), .CK(clk), .Q(instr[23]) );
  DFF_X1 instr_reg_22_ ( .D(in[22]), .CK(clk), .Q(instr[22]) );
  DFF_X1 instr_reg_21_ ( .D(in[21]), .CK(clk), .Q(instr[21]) );
  DFF_X1 instr_reg_20_ ( .D(in[20]), .CK(clk), .Q(instr[20]) );
  DFF_X1 instr_reg_19_ ( .D(in[19]), .CK(clk), .Q(instr[19]) );
  DFF_X1 instr_reg_18_ ( .D(in[18]), .CK(clk), .Q(instr[18]) );
  DFF_X1 instr_reg_17_ ( .D(in[17]), .CK(clk), .Q(instr[17]) );
  DFF_X1 instr_reg_16_ ( .D(in[16]), .CK(clk), .Q(instr[16]) );
  DFF_X1 instr_reg_15_ ( .D(in[15]), .CK(clk), .Q(instr[15]) );
  DFF_X1 instr_reg_14_ ( .D(in[14]), .CK(clk), .Q(instr[14]) );
  DFF_X1 instr_reg_13_ ( .D(in[13]), .CK(clk), .Q(instr[13]) );
  DFF_X1 instr_reg_12_ ( .D(in[12]), .CK(clk), .Q(instr[12]) );
  DFF_X1 instr_reg_11_ ( .D(in[11]), .CK(clk), .Q(instr[11]) );
  DFF_X1 instr_reg_10_ ( .D(in[10]), .CK(clk), .Q(instr[10]) );
  DFF_X1 instr_reg_9_ ( .D(in[9]), .CK(clk), .Q(instr[9]) );
  DFF_X1 instr_reg_8_ ( .D(in[8]), .CK(clk), .Q(instr[8]) );
  DFF_X1 instr_reg_7_ ( .D(in[7]), .CK(clk), .Q(instr[7]) );
  DFF_X1 instr_reg_6_ ( .D(in[6]), .CK(clk), .Q(instr[6]) );
  DFF_X1 instr_reg_5_ ( .D(in[5]), .CK(clk), .Q(instr[5]) );
  DFF_X1 instr_reg_4_ ( .D(in[4]), .CK(clk), .Q(instr[4]) );
  DFF_X1 instr_reg_3_ ( .D(in[3]), .CK(clk), .Q(instr[3]) );
  DFF_X1 instr_reg_2_ ( .D(in[2]), .CK(clk), .Q(instr[2]) );
  DFF_X1 instr_reg_1_ ( .D(in[1]), .CK(clk), .Q(instr[1]) );
  DFF_X1 instr_reg_0_ ( .D(in[0]), .CK(clk), .Q(instr[0]) );
endmodule


module regfile ( clk, ra1, ra2, en_write, wa, wdata, rd1, rd2 );
  input [4:0] ra1;
  input [4:0] ra2;
  input [4:0] wa;
  input [31:0] wdata;
  output [31:0] rd1;
  output [31:0] rd2;
  input clk, en_write;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2286, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2359, n2360, n2362,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2500, n2501, n2503, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2642, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n90, n91, n99, n100, n108, n109, n117, n118, n126, n127, n135, n136,
         n144, n145, n153, n154, n162, n163, n171, n172, n180, n181, n189,
         n190, n326, n327, n335, n336, n344, n345, n353, n354, n362, n363,
         n371, n372, n380, n381, n389, n390, n398, n399, n407, n408, n416,
         n417, n425, n426, n434, n435, n443, n444, n580, n581, n589, n590,
         n598, n599, n607, n608, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n2285,
         n2287, n2357, n2358, n2361, n2363, n2498, n2499, n2502, n2504, n2639,
         n2640, n2641, n2643, n2777, n2778, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724;
  wire   [31:0] x1_ra_w;
  wire   [31:0] x6_t1_w;
  wire   [31:0] x7_t2_w;
  wire   [31:0] x8_s0_w;
  wire   [31:0] x9_s1_w;
  wire   [31:0] x14_a4_w;
  wire   [31:0] x15_a5_w;
  wire   [31:0] x16_a6_w;
  wire   [31:0] x17_a7_w;
  wire   [31:0] x22_s6_w;
  wire   [31:0] x23_s7_w;
  wire   [31:0] x26_s10_w;
  wire   [31:0] x27_s11_w;
  wire   [31:0] x30_t5_w;
  wire   [31:0] x31_t6_w;

  DFF_X1 reg_r28_q_reg_31_ ( .D(n3290), .CK(n3724), .QN(n1) );
  DFF_X1 reg_r28_q_reg_30_ ( .D(n3289), .CK(n3724), .QN(n2) );
  DFF_X1 reg_r28_q_reg_29_ ( .D(n3288), .CK(n3724), .QN(n3) );
  DFF_X1 reg_r28_q_reg_28_ ( .D(n3287), .CK(n3724), .QN(n4) );
  DFF_X1 reg_r28_q_reg_27_ ( .D(n3286), .CK(n3724), .QN(n5) );
  DFF_X1 reg_r28_q_reg_26_ ( .D(n3285), .CK(n3724), .QN(n6) );
  DFF_X1 reg_r28_q_reg_25_ ( .D(n3284), .CK(n3724), .QN(n7) );
  DFF_X1 reg_r28_q_reg_24_ ( .D(n3283), .CK(n3724), .QN(n8) );
  DFF_X1 reg_r28_q_reg_23_ ( .D(n3282), .CK(n3724), .QN(n9) );
  DFF_X1 reg_r28_q_reg_22_ ( .D(n3281), .CK(n3724), .QN(n10) );
  DFF_X1 reg_r28_q_reg_21_ ( .D(n3280), .CK(n3724), .QN(n11) );
  DFF_X1 reg_r28_q_reg_20_ ( .D(n3279), .CK(n3724), .QN(n12) );
  DFF_X1 reg_r28_q_reg_19_ ( .D(n3278), .CK(n3724), .QN(n13) );
  DFF_X1 reg_r28_q_reg_18_ ( .D(n3277), .CK(n3724), .QN(n14) );
  DFF_X1 reg_r28_q_reg_17_ ( .D(n3276), .CK(n3724), .QN(n15) );
  DFF_X1 reg_r28_q_reg_16_ ( .D(n3275), .CK(n3724), .QN(n16) );
  DFF_X1 reg_r28_q_reg_15_ ( .D(n3274), .CK(n3724), .QN(n17) );
  DFF_X1 reg_r28_q_reg_14_ ( .D(n3273), .CK(n3724), .QN(n18) );
  DFF_X1 reg_r28_q_reg_13_ ( .D(n3272), .CK(n3724), .QN(n19) );
  DFF_X1 reg_r28_q_reg_12_ ( .D(n3271), .CK(n3724), .QN(n20) );
  DFF_X1 reg_r28_q_reg_11_ ( .D(n3270), .CK(n3724), .QN(n21) );
  DFF_X1 reg_r28_q_reg_10_ ( .D(n3269), .CK(n3724), .QN(n22) );
  DFF_X1 reg_r28_q_reg_9_ ( .D(n3268), .CK(n3724), .QN(n23) );
  DFF_X1 reg_r28_q_reg_8_ ( .D(n3267), .CK(n3724), .QN(n24) );
  DFF_X1 reg_r28_q_reg_7_ ( .D(n3266), .CK(n3724), .QN(n25) );
  DFF_X1 reg_r28_q_reg_6_ ( .D(n3265), .CK(n3724), .QN(n26) );
  DFF_X1 reg_r28_q_reg_5_ ( .D(n3264), .CK(n3724), .QN(n27) );
  DFF_X1 reg_r28_q_reg_4_ ( .D(n3263), .CK(n3724), .QN(n28) );
  DFF_X1 reg_r28_q_reg_3_ ( .D(n3262), .CK(n3724), .QN(n29) );
  DFF_X1 reg_r28_q_reg_2_ ( .D(n3261), .CK(n3724), .QN(n30) );
  DFF_X1 reg_r28_q_reg_1_ ( .D(n3260), .CK(n3724), .QN(n31) );
  DFF_X1 reg_r28_q_reg_0_ ( .D(n3259), .CK(n3724), .QN(n32) );
  DFF_X1 reg_r29_q_reg_31_ ( .D(n3258), .CK(n3724), .QN(n33) );
  DFF_X1 reg_r29_q_reg_30_ ( .D(n3257), .CK(n3724), .QN(n34) );
  DFF_X1 reg_r29_q_reg_29_ ( .D(n3256), .CK(n3724), .QN(n35) );
  DFF_X1 reg_r29_q_reg_28_ ( .D(n3255), .CK(n3724), .QN(n36) );
  DFF_X1 reg_r29_q_reg_27_ ( .D(n3254), .CK(n3724), .QN(n37) );
  DFF_X1 reg_r29_q_reg_26_ ( .D(n3253), .CK(n3724), .QN(n38) );
  DFF_X1 reg_r29_q_reg_25_ ( .D(n3252), .CK(n3724), .QN(n39) );
  DFF_X1 reg_r29_q_reg_24_ ( .D(n3251), .CK(n3724), .QN(n40) );
  DFF_X1 reg_r29_q_reg_23_ ( .D(n3250), .CK(n3724), .QN(n41) );
  DFF_X1 reg_r29_q_reg_22_ ( .D(n3249), .CK(n3724), .QN(n42) );
  DFF_X1 reg_r29_q_reg_21_ ( .D(n3248), .CK(n3724), .QN(n43) );
  DFF_X1 reg_r29_q_reg_20_ ( .D(n3247), .CK(n3724), .QN(n44) );
  DFF_X1 reg_r29_q_reg_19_ ( .D(n3246), .CK(n3724), .QN(n45) );
  DFF_X1 reg_r29_q_reg_18_ ( .D(n3245), .CK(n3724), .QN(n46) );
  DFF_X1 reg_r29_q_reg_17_ ( .D(n3244), .CK(n3724), .QN(n47) );
  DFF_X1 reg_r29_q_reg_16_ ( .D(n3243), .CK(n3724), .QN(n48) );
  DFF_X1 reg_r29_q_reg_15_ ( .D(n3242), .CK(n3724), .QN(n49) );
  DFF_X1 reg_r29_q_reg_14_ ( .D(n3241), .CK(n3724), .QN(n50) );
  DFF_X1 reg_r29_q_reg_13_ ( .D(n3240), .CK(n3724), .QN(n51) );
  DFF_X1 reg_r29_q_reg_12_ ( .D(n3239), .CK(n3724), .QN(n52) );
  DFF_X1 reg_r29_q_reg_11_ ( .D(n3238), .CK(n3724), .QN(n53) );
  DFF_X1 reg_r29_q_reg_10_ ( .D(n3237), .CK(n3724), .QN(n54) );
  DFF_X1 reg_r29_q_reg_9_ ( .D(n3236), .CK(n3724), .QN(n55) );
  DFF_X1 reg_r29_q_reg_8_ ( .D(n3235), .CK(n3724), .QN(n56) );
  DFF_X1 reg_r29_q_reg_7_ ( .D(n3234), .CK(n3724), .QN(n57) );
  DFF_X1 reg_r29_q_reg_6_ ( .D(n3233), .CK(n3724), .QN(n58) );
  DFF_X1 reg_r29_q_reg_5_ ( .D(n3232), .CK(n3724), .QN(n59) );
  DFF_X1 reg_r29_q_reg_4_ ( .D(n3231), .CK(n3724), .QN(n60) );
  DFF_X1 reg_r29_q_reg_3_ ( .D(n3230), .CK(n3724), .QN(n61) );
  DFF_X1 reg_r29_q_reg_2_ ( .D(n3229), .CK(n3724), .QN(n62) );
  DFF_X1 reg_r29_q_reg_1_ ( .D(n3228), .CK(n3724), .QN(n63) );
  DFF_X1 reg_r29_q_reg_0_ ( .D(n3227), .CK(n3724), .QN(n64) );
  DFF_X1 reg_r27_q_reg_31_ ( .D(n995), .CK(n3724), .Q(x27_s11_w[31]) );
  DFF_X1 reg_r27_q_reg_30_ ( .D(n1011), .CK(n3724), .Q(x27_s11_w[30]) );
  DFF_X1 reg_r27_q_reg_29_ ( .D(n1027), .CK(n3724), .Q(x27_s11_w[29]) );
  DFF_X1 reg_r27_q_reg_28_ ( .D(n1043), .CK(n3724), .Q(x27_s11_w[28]) );
  DFF_X1 reg_r27_q_reg_27_ ( .D(n1059), .CK(n3724), .Q(x27_s11_w[27]) );
  DFF_X1 reg_r27_q_reg_26_ ( .D(n2363), .CK(n3724), .Q(x27_s11_w[26]) );
  DFF_X1 reg_r27_q_reg_25_ ( .D(n3296), .CK(n3724), .Q(x27_s11_w[25]) );
  DFF_X1 reg_r27_q_reg_24_ ( .D(n3312), .CK(n3724), .Q(x27_s11_w[24]) );
  DFF_X1 reg_r27_q_reg_23_ ( .D(n3328), .CK(n3724), .Q(x27_s11_w[23]) );
  DFF_X1 reg_r27_q_reg_22_ ( .D(n3344), .CK(n3724), .Q(x27_s11_w[22]) );
  DFF_X1 reg_r27_q_reg_21_ ( .D(n3360), .CK(n3724), .Q(x27_s11_w[21]) );
  DFF_X1 reg_r27_q_reg_20_ ( .D(n3376), .CK(n3724), .Q(x27_s11_w[20]) );
  DFF_X1 reg_r27_q_reg_19_ ( .D(n3392), .CK(n3724), .Q(x27_s11_w[19]) );
  DFF_X1 reg_r27_q_reg_18_ ( .D(n3408), .CK(n3724), .Q(x27_s11_w[18]) );
  DFF_X1 reg_r27_q_reg_17_ ( .D(n3424), .CK(n3724), .Q(x27_s11_w[17]) );
  DFF_X1 reg_r27_q_reg_16_ ( .D(n3440), .CK(n3724), .Q(x27_s11_w[16]) );
  DFF_X1 reg_r27_q_reg_15_ ( .D(n3456), .CK(n3724), .Q(x27_s11_w[15]) );
  DFF_X1 reg_r27_q_reg_14_ ( .D(n3472), .CK(n3724), .Q(x27_s11_w[14]) );
  DFF_X1 reg_r27_q_reg_13_ ( .D(n3488), .CK(n3724), .Q(x27_s11_w[13]) );
  DFF_X1 reg_r27_q_reg_12_ ( .D(n3504), .CK(n3724), .Q(x27_s11_w[12]) );
  DFF_X1 reg_r27_q_reg_11_ ( .D(n3520), .CK(n3724), .Q(x27_s11_w[11]) );
  DFF_X1 reg_r27_q_reg_10_ ( .D(n3536), .CK(n3724), .Q(x27_s11_w[10]) );
  DFF_X1 reg_r27_q_reg_9_ ( .D(n3552), .CK(n3724), .Q(x27_s11_w[9]) );
  DFF_X1 reg_r27_q_reg_8_ ( .D(n3568), .CK(n3724), .Q(x27_s11_w[8]) );
  DFF_X1 reg_r27_q_reg_7_ ( .D(n3584), .CK(n3724), .Q(x27_s11_w[7]) );
  DFF_X1 reg_r27_q_reg_6_ ( .D(n3600), .CK(n3724), .Q(x27_s11_w[6]) );
  DFF_X1 reg_r27_q_reg_5_ ( .D(n3616), .CK(n3724), .Q(x27_s11_w[5]) );
  DFF_X1 reg_r27_q_reg_4_ ( .D(n3632), .CK(n3724), .Q(x27_s11_w[4]) );
  DFF_X1 reg_r27_q_reg_3_ ( .D(n3648), .CK(n3724), .Q(x27_s11_w[3]) );
  DFF_X1 reg_r27_q_reg_2_ ( .D(n3664), .CK(n3724), .Q(x27_s11_w[2]) );
  DFF_X1 reg_r27_q_reg_1_ ( .D(n3680), .CK(n3724), .Q(x27_s11_w[1]) );
  DFF_X1 reg_r27_q_reg_0_ ( .D(n3696), .CK(n3724), .Q(x27_s11_w[0]) );
  DFF_X1 reg_r30_q_reg_31_ ( .D(n996), .CK(n3724), .Q(x30_t5_w[31]) );
  DFF_X1 reg_r30_q_reg_30_ ( .D(n1012), .CK(n3724), .Q(x30_t5_w[30]) );
  DFF_X1 reg_r30_q_reg_29_ ( .D(n1028), .CK(n3724), .Q(x30_t5_w[29]) );
  DFF_X1 reg_r30_q_reg_28_ ( .D(n1044), .CK(n3724), .Q(x30_t5_w[28]) );
  DFF_X1 reg_r30_q_reg_27_ ( .D(n1060), .CK(n3724), .Q(x30_t5_w[27]) );
  DFF_X1 reg_r30_q_reg_26_ ( .D(n2498), .CK(n3724), .Q(x30_t5_w[26]) );
  DFF_X1 reg_r30_q_reg_25_ ( .D(n3297), .CK(n3724), .Q(x30_t5_w[25]) );
  DFF_X1 reg_r30_q_reg_24_ ( .D(n3313), .CK(n3724), .Q(x30_t5_w[24]) );
  DFF_X1 reg_r30_q_reg_23_ ( .D(n3329), .CK(n3724), .Q(x30_t5_w[23]) );
  DFF_X1 reg_r30_q_reg_22_ ( .D(n3345), .CK(n3724), .Q(x30_t5_w[22]) );
  DFF_X1 reg_r30_q_reg_21_ ( .D(n3361), .CK(n3724), .Q(x30_t5_w[21]) );
  DFF_X1 reg_r30_q_reg_20_ ( .D(n3377), .CK(n3724), .Q(x30_t5_w[20]) );
  DFF_X1 reg_r30_q_reg_19_ ( .D(n3393), .CK(n3724), .Q(x30_t5_w[19]) );
  DFF_X1 reg_r30_q_reg_18_ ( .D(n3409), .CK(n3724), .Q(x30_t5_w[18]) );
  DFF_X1 reg_r30_q_reg_17_ ( .D(n3425), .CK(n3724), .Q(x30_t5_w[17]) );
  DFF_X1 reg_r30_q_reg_16_ ( .D(n3441), .CK(n3724), .Q(x30_t5_w[16]) );
  DFF_X1 reg_r30_q_reg_15_ ( .D(n3457), .CK(n3724), .Q(x30_t5_w[15]) );
  DFF_X1 reg_r30_q_reg_14_ ( .D(n3473), .CK(n3724), .Q(x30_t5_w[14]) );
  DFF_X1 reg_r30_q_reg_13_ ( .D(n3489), .CK(n3724), .Q(x30_t5_w[13]) );
  DFF_X1 reg_r30_q_reg_12_ ( .D(n3505), .CK(n3724), .Q(x30_t5_w[12]) );
  DFF_X1 reg_r30_q_reg_11_ ( .D(n3521), .CK(n3724), .Q(x30_t5_w[11]) );
  DFF_X1 reg_r30_q_reg_10_ ( .D(n3537), .CK(n3724), .Q(x30_t5_w[10]) );
  DFF_X1 reg_r30_q_reg_9_ ( .D(n3553), .CK(n3724), .Q(x30_t5_w[9]) );
  DFF_X1 reg_r30_q_reg_8_ ( .D(n3569), .CK(n3724), .Q(x30_t5_w[8]) );
  DFF_X1 reg_r30_q_reg_7_ ( .D(n3585), .CK(n3724), .Q(x30_t5_w[7]) );
  DFF_X1 reg_r30_q_reg_6_ ( .D(n3601), .CK(n3724), .Q(x30_t5_w[6]) );
  DFF_X1 reg_r30_q_reg_5_ ( .D(n3617), .CK(n3724), .Q(x30_t5_w[5]) );
  DFF_X1 reg_r30_q_reg_4_ ( .D(n3633), .CK(n3724), .Q(x30_t5_w[4]) );
  DFF_X1 reg_r30_q_reg_3_ ( .D(n3649), .CK(n3724), .Q(x30_t5_w[3]) );
  DFF_X1 reg_r30_q_reg_2_ ( .D(n3665), .CK(n3724), .Q(x30_t5_w[2]) );
  DFF_X1 reg_r30_q_reg_1_ ( .D(n3681), .CK(n3724), .Q(x30_t5_w[1]) );
  DFF_X1 reg_r30_q_reg_0_ ( .D(n3697), .CK(n3724), .Q(x30_t5_w[0]) );
  DFF_X1 reg_r31_q_reg_31_ ( .D(n997), .CK(n3724), .Q(x31_t6_w[31]) );
  DFF_X1 reg_r31_q_reg_30_ ( .D(n1013), .CK(n3724), .Q(x31_t6_w[30]) );
  DFF_X1 reg_r31_q_reg_29_ ( .D(n1029), .CK(n3724), .Q(x31_t6_w[29]) );
  DFF_X1 reg_r31_q_reg_28_ ( .D(n1045), .CK(n3724), .Q(x31_t6_w[28]) );
  DFF_X1 reg_r31_q_reg_27_ ( .D(n1061), .CK(n3724), .Q(x31_t6_w[27]) );
  DFF_X1 reg_r31_q_reg_26_ ( .D(n2499), .CK(n3724), .Q(x31_t6_w[26]) );
  DFF_X1 reg_r31_q_reg_25_ ( .D(n3298), .CK(n3724), .Q(x31_t6_w[25]) );
  DFF_X1 reg_r31_q_reg_24_ ( .D(n3314), .CK(n3724), .Q(x31_t6_w[24]) );
  DFF_X1 reg_r31_q_reg_23_ ( .D(n3330), .CK(n3724), .Q(x31_t6_w[23]) );
  DFF_X1 reg_r31_q_reg_22_ ( .D(n3346), .CK(n3724), .Q(x31_t6_w[22]) );
  DFF_X1 reg_r31_q_reg_21_ ( .D(n3362), .CK(n3724), .Q(x31_t6_w[21]) );
  DFF_X1 reg_r31_q_reg_20_ ( .D(n3378), .CK(n3724), .Q(x31_t6_w[20]) );
  DFF_X1 reg_r31_q_reg_19_ ( .D(n3394), .CK(n3724), .Q(x31_t6_w[19]) );
  DFF_X1 reg_r31_q_reg_18_ ( .D(n3410), .CK(n3724), .Q(x31_t6_w[18]) );
  DFF_X1 reg_r31_q_reg_17_ ( .D(n3426), .CK(n3724), .Q(x31_t6_w[17]) );
  DFF_X1 reg_r31_q_reg_16_ ( .D(n3442), .CK(n3724), .Q(x31_t6_w[16]) );
  DFF_X1 reg_r31_q_reg_15_ ( .D(n3458), .CK(n3724), .Q(x31_t6_w[15]) );
  DFF_X1 reg_r31_q_reg_14_ ( .D(n3474), .CK(n3724), .Q(x31_t6_w[14]) );
  DFF_X1 reg_r31_q_reg_13_ ( .D(n3490), .CK(n3724), .Q(x31_t6_w[13]) );
  DFF_X1 reg_r31_q_reg_12_ ( .D(n3506), .CK(n3724), .Q(x31_t6_w[12]) );
  DFF_X1 reg_r31_q_reg_11_ ( .D(n3522), .CK(n3724), .Q(x31_t6_w[11]) );
  DFF_X1 reg_r31_q_reg_10_ ( .D(n3538), .CK(n3724), .Q(x31_t6_w[10]) );
  DFF_X1 reg_r31_q_reg_9_ ( .D(n3554), .CK(n3724), .Q(x31_t6_w[9]) );
  DFF_X1 reg_r31_q_reg_8_ ( .D(n3570), .CK(n3724), .Q(x31_t6_w[8]) );
  DFF_X1 reg_r31_q_reg_7_ ( .D(n3586), .CK(n3724), .Q(x31_t6_w[7]) );
  DFF_X1 reg_r31_q_reg_6_ ( .D(n3602), .CK(n3724), .Q(x31_t6_w[6]) );
  DFF_X1 reg_r31_q_reg_5_ ( .D(n3618), .CK(n3724), .Q(x31_t6_w[5]) );
  DFF_X1 reg_r31_q_reg_4_ ( .D(n3634), .CK(n3724), .Q(x31_t6_w[4]) );
  DFF_X1 reg_r31_q_reg_3_ ( .D(n3650), .CK(n3724), .Q(x31_t6_w[3]) );
  DFF_X1 reg_r31_q_reg_2_ ( .D(n3666), .CK(n3724), .Q(x31_t6_w[2]) );
  DFF_X1 reg_r31_q_reg_1_ ( .D(n3682), .CK(n3724), .Q(x31_t6_w[1]) );
  DFF_X1 reg_r31_q_reg_0_ ( .D(n3698), .CK(n3724), .Q(x31_t6_w[0]) );
  DFF_X1 reg_r1_q_reg_31_ ( .D(n998), .CK(n3724), .Q(x1_ra_w[31]) );
  DFF_X1 reg_r1_q_reg_30_ ( .D(n1014), .CK(n3724), .Q(x1_ra_w[30]) );
  DFF_X1 reg_r1_q_reg_29_ ( .D(n1030), .CK(n3724), .Q(x1_ra_w[29]) );
  DFF_X1 reg_r1_q_reg_28_ ( .D(n1046), .CK(n3724), .Q(x1_ra_w[28]) );
  DFF_X1 reg_r1_q_reg_27_ ( .D(n1062), .CK(n3724), .Q(x1_ra_w[27]) );
  DFF_X1 reg_r1_q_reg_26_ ( .D(n2502), .CK(n3724), .Q(x1_ra_w[26]) );
  DFF_X1 reg_r1_q_reg_25_ ( .D(n3299), .CK(n3724), .Q(x1_ra_w[25]) );
  DFF_X1 reg_r1_q_reg_24_ ( .D(n3315), .CK(n3724), .Q(x1_ra_w[24]) );
  DFF_X1 reg_r1_q_reg_23_ ( .D(n3331), .CK(n3724), .Q(x1_ra_w[23]) );
  DFF_X1 reg_r1_q_reg_22_ ( .D(n3347), .CK(n3724), .Q(x1_ra_w[22]) );
  DFF_X1 reg_r1_q_reg_21_ ( .D(n3363), .CK(n3724), .Q(x1_ra_w[21]) );
  DFF_X1 reg_r1_q_reg_20_ ( .D(n3379), .CK(n3724), .Q(x1_ra_w[20]) );
  DFF_X1 reg_r1_q_reg_19_ ( .D(n3395), .CK(n3724), .Q(x1_ra_w[19]) );
  DFF_X1 reg_r1_q_reg_18_ ( .D(n3411), .CK(n3724), .Q(x1_ra_w[18]) );
  DFF_X1 reg_r1_q_reg_17_ ( .D(n3427), .CK(n3724), .Q(x1_ra_w[17]) );
  DFF_X1 reg_r1_q_reg_16_ ( .D(n3443), .CK(n3724), .Q(x1_ra_w[16]) );
  DFF_X1 reg_r1_q_reg_15_ ( .D(n3459), .CK(n3724), .Q(x1_ra_w[15]) );
  DFF_X1 reg_r1_q_reg_14_ ( .D(n3475), .CK(n3724), .Q(x1_ra_w[14]) );
  DFF_X1 reg_r1_q_reg_13_ ( .D(n3491), .CK(n3724), .Q(x1_ra_w[13]) );
  DFF_X1 reg_r1_q_reg_12_ ( .D(n3507), .CK(n3724), .Q(x1_ra_w[12]) );
  DFF_X1 reg_r1_q_reg_11_ ( .D(n3523), .CK(n3724), .Q(x1_ra_w[11]) );
  DFF_X1 reg_r1_q_reg_10_ ( .D(n3539), .CK(n3724), .Q(x1_ra_w[10]) );
  DFF_X1 reg_r1_q_reg_9_ ( .D(n3555), .CK(n3724), .Q(x1_ra_w[9]) );
  DFF_X1 reg_r1_q_reg_8_ ( .D(n3571), .CK(n3724), .Q(x1_ra_w[8]) );
  DFF_X1 reg_r1_q_reg_7_ ( .D(n3587), .CK(n3724), .Q(x1_ra_w[7]) );
  DFF_X1 reg_r1_q_reg_6_ ( .D(n3603), .CK(n3724), .Q(x1_ra_w[6]) );
  DFF_X1 reg_r1_q_reg_5_ ( .D(n3619), .CK(n3724), .Q(x1_ra_w[5]) );
  DFF_X1 reg_r1_q_reg_4_ ( .D(n3635), .CK(n3724), .Q(x1_ra_w[4]) );
  DFF_X1 reg_r1_q_reg_3_ ( .D(n3651), .CK(n3724), .Q(x1_ra_w[3]) );
  DFF_X1 reg_r1_q_reg_2_ ( .D(n3667), .CK(n3724), .Q(x1_ra_w[2]) );
  DFF_X1 reg_r1_q_reg_1_ ( .D(n3683), .CK(n3724), .Q(x1_ra_w[1]) );
  DFF_X1 reg_r1_q_reg_0_ ( .D(n3699), .CK(n3724), .Q(x1_ra_w[0]) );
  DFF_X1 reg_r2_q_reg_31_ ( .D(n3226), .CK(n3724), .QN(n193) );
  DFF_X1 reg_r2_q_reg_30_ ( .D(n3225), .CK(n3724), .QN(n194) );
  DFF_X1 reg_r2_q_reg_29_ ( .D(n3224), .CK(n3724), .QN(n195) );
  DFF_X1 reg_r2_q_reg_28_ ( .D(n3223), .CK(n3724), .QN(n196) );
  DFF_X1 reg_r2_q_reg_27_ ( .D(n3222), .CK(n3724), .QN(n197) );
  DFF_X1 reg_r2_q_reg_26_ ( .D(n3221), .CK(n3724), .QN(n198) );
  DFF_X1 reg_r2_q_reg_25_ ( .D(n3220), .CK(n3724), .QN(n199) );
  DFF_X1 reg_r2_q_reg_24_ ( .D(n3219), .CK(n3724), .QN(n200) );
  DFF_X1 reg_r2_q_reg_23_ ( .D(n3218), .CK(n3724), .QN(n201) );
  DFF_X1 reg_r2_q_reg_22_ ( .D(n3217), .CK(n3724), .QN(n202) );
  DFF_X1 reg_r2_q_reg_21_ ( .D(n3216), .CK(n3724), .QN(n203) );
  DFF_X1 reg_r2_q_reg_20_ ( .D(n3215), .CK(n3724), .QN(n204) );
  DFF_X1 reg_r2_q_reg_19_ ( .D(n3214), .CK(n3724), .QN(n205) );
  DFF_X1 reg_r2_q_reg_18_ ( .D(n3213), .CK(n3724), .QN(n206) );
  DFF_X1 reg_r2_q_reg_17_ ( .D(n3212), .CK(n3724), .QN(n207) );
  DFF_X1 reg_r2_q_reg_16_ ( .D(n3211), .CK(n3724), .QN(n208) );
  DFF_X1 reg_r2_q_reg_15_ ( .D(n3210), .CK(n3724), .QN(n209) );
  DFF_X1 reg_r2_q_reg_14_ ( .D(n3209), .CK(n3724), .QN(n210) );
  DFF_X1 reg_r2_q_reg_13_ ( .D(n3208), .CK(n3724), .QN(n211) );
  DFF_X1 reg_r2_q_reg_12_ ( .D(n3207), .CK(n3724), .QN(n212) );
  DFF_X1 reg_r2_q_reg_11_ ( .D(n3206), .CK(n3724), .QN(n213) );
  DFF_X1 reg_r2_q_reg_10_ ( .D(n3205), .CK(n3724), .QN(n214) );
  DFF_X1 reg_r2_q_reg_9_ ( .D(n3204), .CK(n3724), .QN(n215) );
  DFF_X1 reg_r2_q_reg_8_ ( .D(n3203), .CK(n3724), .QN(n216) );
  DFF_X1 reg_r2_q_reg_7_ ( .D(n3202), .CK(n3724), .QN(n217) );
  DFF_X1 reg_r2_q_reg_6_ ( .D(n3201), .CK(n3724), .QN(n218) );
  DFF_X1 reg_r2_q_reg_5_ ( .D(n3200), .CK(n3724), .QN(n219) );
  DFF_X1 reg_r2_q_reg_4_ ( .D(n3199), .CK(n3724), .QN(n220) );
  DFF_X1 reg_r2_q_reg_3_ ( .D(n3198), .CK(n3724), .QN(n221) );
  DFF_X1 reg_r2_q_reg_2_ ( .D(n3197), .CK(n3724), .QN(n222) );
  DFF_X1 reg_r2_q_reg_1_ ( .D(n3196), .CK(n3724), .QN(n223) );
  DFF_X1 reg_r2_q_reg_0_ ( .D(n3195), .CK(n3724), .QN(n224) );
  DFF_X1 reg_r3_q_reg_31_ ( .D(n3194), .CK(n3724), .QN(n225) );
  DFF_X1 reg_r3_q_reg_30_ ( .D(n3193), .CK(n3724), .QN(n226) );
  DFF_X1 reg_r3_q_reg_29_ ( .D(n3192), .CK(n3724), .QN(n227) );
  DFF_X1 reg_r3_q_reg_28_ ( .D(n3191), .CK(n3724), .QN(n228) );
  DFF_X1 reg_r3_q_reg_27_ ( .D(n3190), .CK(n3724), .QN(n229) );
  DFF_X1 reg_r3_q_reg_26_ ( .D(n3189), .CK(n3724), .QN(n230) );
  DFF_X1 reg_r3_q_reg_25_ ( .D(n3188), .CK(n3724), .QN(n231) );
  DFF_X1 reg_r3_q_reg_24_ ( .D(n3187), .CK(n3724), .QN(n232) );
  DFF_X1 reg_r3_q_reg_23_ ( .D(n3186), .CK(n3724), .QN(n233) );
  DFF_X1 reg_r3_q_reg_22_ ( .D(n3185), .CK(n3724), .QN(n234) );
  DFF_X1 reg_r3_q_reg_21_ ( .D(n3184), .CK(n3724), .QN(n235) );
  DFF_X1 reg_r3_q_reg_20_ ( .D(n3183), .CK(n3724), .QN(n236) );
  DFF_X1 reg_r3_q_reg_19_ ( .D(n3182), .CK(n3724), .QN(n237) );
  DFF_X1 reg_r3_q_reg_18_ ( .D(n3181), .CK(n3724), .QN(n238) );
  DFF_X1 reg_r3_q_reg_17_ ( .D(n3180), .CK(n3724), .QN(n239) );
  DFF_X1 reg_r3_q_reg_16_ ( .D(n3179), .CK(n3724), .QN(n240) );
  DFF_X1 reg_r3_q_reg_15_ ( .D(n3178), .CK(n3724), .QN(n241) );
  DFF_X1 reg_r3_q_reg_14_ ( .D(n3177), .CK(n3724), .QN(n242) );
  DFF_X1 reg_r3_q_reg_13_ ( .D(n3176), .CK(n3724), .QN(n243) );
  DFF_X1 reg_r3_q_reg_12_ ( .D(n3175), .CK(n3724), .QN(n244) );
  DFF_X1 reg_r3_q_reg_11_ ( .D(n3174), .CK(n3724), .QN(n245) );
  DFF_X1 reg_r3_q_reg_10_ ( .D(n3173), .CK(n3724), .QN(n246) );
  DFF_X1 reg_r3_q_reg_9_ ( .D(n3172), .CK(n3724), .QN(n247) );
  DFF_X1 reg_r3_q_reg_8_ ( .D(n3171), .CK(n3724), .QN(n248) );
  DFF_X1 reg_r3_q_reg_7_ ( .D(n3170), .CK(n3724), .QN(n249) );
  DFF_X1 reg_r3_q_reg_6_ ( .D(n3169), .CK(n3724), .QN(n250) );
  DFF_X1 reg_r3_q_reg_5_ ( .D(n3168), .CK(n3724), .QN(n251) );
  DFF_X1 reg_r3_q_reg_4_ ( .D(n3167), .CK(n3724), .QN(n252) );
  DFF_X1 reg_r3_q_reg_3_ ( .D(n3166), .CK(n3724), .QN(n253) );
  DFF_X1 reg_r3_q_reg_2_ ( .D(n3165), .CK(n3724), .QN(n254) );
  DFF_X1 reg_r3_q_reg_1_ ( .D(n3164), .CK(n3724), .QN(n255) );
  DFF_X1 reg_r3_q_reg_0_ ( .D(n3163), .CK(n3724), .QN(n256) );
  DFF_X1 reg_r4_q_reg_31_ ( .D(n3162), .CK(n3724), .QN(n257) );
  DFF_X1 reg_r4_q_reg_30_ ( .D(n3161), .CK(n3724), .QN(n258) );
  DFF_X1 reg_r4_q_reg_29_ ( .D(n3160), .CK(n3724), .QN(n259) );
  DFF_X1 reg_r4_q_reg_28_ ( .D(n3159), .CK(n3724), .QN(n260) );
  DFF_X1 reg_r4_q_reg_27_ ( .D(n3158), .CK(n3724), .QN(n261) );
  DFF_X1 reg_r4_q_reg_26_ ( .D(n3157), .CK(n3724), .QN(n262) );
  DFF_X1 reg_r4_q_reg_25_ ( .D(n3156), .CK(n3724), .QN(n263) );
  DFF_X1 reg_r4_q_reg_24_ ( .D(n3155), .CK(n3724), .QN(n264) );
  DFF_X1 reg_r4_q_reg_23_ ( .D(n3154), .CK(n3724), .QN(n265) );
  DFF_X1 reg_r4_q_reg_22_ ( .D(n3153), .CK(n3724), .QN(n266) );
  DFF_X1 reg_r4_q_reg_21_ ( .D(n3152), .CK(n3724), .QN(n267) );
  DFF_X1 reg_r4_q_reg_20_ ( .D(n3151), .CK(n3724), .QN(n268) );
  DFF_X1 reg_r4_q_reg_19_ ( .D(n3150), .CK(n3724), .QN(n269) );
  DFF_X1 reg_r4_q_reg_18_ ( .D(n3149), .CK(n3724), .QN(n270) );
  DFF_X1 reg_r4_q_reg_17_ ( .D(n3148), .CK(n3724), .QN(n271) );
  DFF_X1 reg_r4_q_reg_16_ ( .D(n3147), .CK(n3724), .QN(n272) );
  DFF_X1 reg_r4_q_reg_15_ ( .D(n3146), .CK(n3724), .QN(n273) );
  DFF_X1 reg_r4_q_reg_14_ ( .D(n3145), .CK(n3724), .QN(n274) );
  DFF_X1 reg_r4_q_reg_13_ ( .D(n3144), .CK(n3724), .QN(n275) );
  DFF_X1 reg_r4_q_reg_12_ ( .D(n3143), .CK(n3724), .QN(n276) );
  DFF_X1 reg_r4_q_reg_11_ ( .D(n3142), .CK(n3724), .QN(n277) );
  DFF_X1 reg_r4_q_reg_10_ ( .D(n3141), .CK(n3724), .QN(n278) );
  DFF_X1 reg_r4_q_reg_9_ ( .D(n3140), .CK(n3724), .QN(n279) );
  DFF_X1 reg_r4_q_reg_8_ ( .D(n3139), .CK(n3724), .QN(n280) );
  DFF_X1 reg_r4_q_reg_7_ ( .D(n3138), .CK(n3724), .QN(n281) );
  DFF_X1 reg_r4_q_reg_6_ ( .D(n3137), .CK(n3724), .QN(n282) );
  DFF_X1 reg_r4_q_reg_5_ ( .D(n3136), .CK(n3724), .QN(n283) );
  DFF_X1 reg_r4_q_reg_4_ ( .D(n3135), .CK(n3724), .QN(n284) );
  DFF_X1 reg_r4_q_reg_3_ ( .D(n3134), .CK(n3724), .QN(n285) );
  DFF_X1 reg_r4_q_reg_2_ ( .D(n3133), .CK(n3724), .QN(n286) );
  DFF_X1 reg_r4_q_reg_1_ ( .D(n3132), .CK(n3724), .QN(n287) );
  DFF_X1 reg_r4_q_reg_0_ ( .D(n3131), .CK(n3724), .QN(n288) );
  DFF_X1 reg_r5_q_reg_31_ ( .D(n3130), .CK(n3724), .QN(n289) );
  DFF_X1 reg_r5_q_reg_30_ ( .D(n3129), .CK(n3724), .QN(n290) );
  DFF_X1 reg_r5_q_reg_29_ ( .D(n3128), .CK(n3724), .QN(n291) );
  DFF_X1 reg_r5_q_reg_28_ ( .D(n3127), .CK(n3724), .QN(n292) );
  DFF_X1 reg_r5_q_reg_27_ ( .D(n3126), .CK(n3724), .QN(n293) );
  DFF_X1 reg_r5_q_reg_26_ ( .D(n3125), .CK(n3724), .QN(n294) );
  DFF_X1 reg_r5_q_reg_25_ ( .D(n3124), .CK(n3724), .QN(n295) );
  DFF_X1 reg_r5_q_reg_24_ ( .D(n3123), .CK(n3724), .QN(n296) );
  DFF_X1 reg_r5_q_reg_23_ ( .D(n3122), .CK(n3724), .QN(n297) );
  DFF_X1 reg_r5_q_reg_22_ ( .D(n3121), .CK(n3724), .QN(n298) );
  DFF_X1 reg_r5_q_reg_21_ ( .D(n3120), .CK(n3724), .QN(n299) );
  DFF_X1 reg_r5_q_reg_20_ ( .D(n3119), .CK(n3724), .QN(n300) );
  DFF_X1 reg_r5_q_reg_19_ ( .D(n3118), .CK(n3724), .QN(n301) );
  DFF_X1 reg_r5_q_reg_18_ ( .D(n3117), .CK(n3724), .QN(n302) );
  DFF_X1 reg_r5_q_reg_17_ ( .D(n3116), .CK(n3724), .QN(n303) );
  DFF_X1 reg_r5_q_reg_16_ ( .D(n3115), .CK(n3724), .QN(n304) );
  DFF_X1 reg_r5_q_reg_15_ ( .D(n3114), .CK(n3724), .QN(n305) );
  DFF_X1 reg_r5_q_reg_14_ ( .D(n3113), .CK(n3724), .QN(n306) );
  DFF_X1 reg_r5_q_reg_13_ ( .D(n3112), .CK(n3724), .QN(n307) );
  DFF_X1 reg_r5_q_reg_12_ ( .D(n3111), .CK(n3724), .QN(n308) );
  DFF_X1 reg_r5_q_reg_11_ ( .D(n3110), .CK(n3724), .QN(n309) );
  DFF_X1 reg_r5_q_reg_10_ ( .D(n3109), .CK(n3724), .QN(n310) );
  DFF_X1 reg_r5_q_reg_9_ ( .D(n3108), .CK(n3724), .QN(n311) );
  DFF_X1 reg_r5_q_reg_8_ ( .D(n3107), .CK(n3724), .QN(n312) );
  DFF_X1 reg_r5_q_reg_7_ ( .D(n3106), .CK(n3724), .QN(n313) );
  DFF_X1 reg_r5_q_reg_6_ ( .D(n3105), .CK(n3724), .QN(n314) );
  DFF_X1 reg_r5_q_reg_5_ ( .D(n3104), .CK(n3724), .QN(n315) );
  DFF_X1 reg_r5_q_reg_4_ ( .D(n3103), .CK(n3724), .QN(n316) );
  DFF_X1 reg_r5_q_reg_3_ ( .D(n3102), .CK(n3724), .QN(n317) );
  DFF_X1 reg_r5_q_reg_2_ ( .D(n3101), .CK(n3724), .QN(n318) );
  DFF_X1 reg_r5_q_reg_1_ ( .D(n3100), .CK(n3724), .QN(n319) );
  DFF_X1 reg_r5_q_reg_0_ ( .D(n3099), .CK(n3724), .QN(n320) );
  DFF_X1 reg_r6_q_reg_31_ ( .D(n999), .CK(n3724), .Q(x6_t1_w[31]) );
  DFF_X1 reg_r6_q_reg_30_ ( .D(n1015), .CK(n3724), .Q(x6_t1_w[30]) );
  DFF_X1 reg_r6_q_reg_29_ ( .D(n1031), .CK(n3724), .Q(x6_t1_w[29]) );
  DFF_X1 reg_r6_q_reg_28_ ( .D(n1047), .CK(n3724), .Q(x6_t1_w[28]) );
  DFF_X1 reg_r6_q_reg_27_ ( .D(n1063), .CK(n3724), .Q(x6_t1_w[27]) );
  DFF_X1 reg_r6_q_reg_26_ ( .D(n2504), .CK(n3724), .Q(x6_t1_w[26]) );
  DFF_X1 reg_r6_q_reg_25_ ( .D(n3300), .CK(n3724), .Q(x6_t1_w[25]) );
  DFF_X1 reg_r6_q_reg_24_ ( .D(n3316), .CK(n3724), .Q(x6_t1_w[24]) );
  DFF_X1 reg_r6_q_reg_23_ ( .D(n3332), .CK(n3724), .Q(x6_t1_w[23]) );
  DFF_X1 reg_r6_q_reg_22_ ( .D(n3348), .CK(n3724), .Q(x6_t1_w[22]) );
  DFF_X1 reg_r6_q_reg_21_ ( .D(n3364), .CK(n3724), .Q(x6_t1_w[21]) );
  DFF_X1 reg_r6_q_reg_20_ ( .D(n3380), .CK(n3724), .Q(x6_t1_w[20]) );
  DFF_X1 reg_r6_q_reg_19_ ( .D(n3396), .CK(n3724), .Q(x6_t1_w[19]) );
  DFF_X1 reg_r6_q_reg_18_ ( .D(n3412), .CK(n3724), .Q(x6_t1_w[18]) );
  DFF_X1 reg_r6_q_reg_17_ ( .D(n3428), .CK(n3724), .Q(x6_t1_w[17]) );
  DFF_X1 reg_r6_q_reg_16_ ( .D(n3444), .CK(n3724), .Q(x6_t1_w[16]) );
  DFF_X1 reg_r6_q_reg_15_ ( .D(n3460), .CK(n3724), .Q(x6_t1_w[15]) );
  DFF_X1 reg_r6_q_reg_14_ ( .D(n3476), .CK(n3724), .Q(x6_t1_w[14]) );
  DFF_X1 reg_r6_q_reg_13_ ( .D(n3492), .CK(n3724), .Q(x6_t1_w[13]) );
  DFF_X1 reg_r6_q_reg_12_ ( .D(n3508), .CK(n3724), .Q(x6_t1_w[12]) );
  DFF_X1 reg_r6_q_reg_11_ ( .D(n3524), .CK(n3724), .Q(x6_t1_w[11]) );
  DFF_X1 reg_r6_q_reg_10_ ( .D(n3540), .CK(n3724), .Q(x6_t1_w[10]) );
  DFF_X1 reg_r6_q_reg_9_ ( .D(n3556), .CK(n3724), .Q(x6_t1_w[9]) );
  DFF_X1 reg_r6_q_reg_8_ ( .D(n3572), .CK(n3724), .Q(x6_t1_w[8]) );
  DFF_X1 reg_r6_q_reg_7_ ( .D(n3588), .CK(n3724), .Q(x6_t1_w[7]) );
  DFF_X1 reg_r6_q_reg_6_ ( .D(n3604), .CK(n3724), .Q(x6_t1_w[6]) );
  DFF_X1 reg_r6_q_reg_5_ ( .D(n3620), .CK(n3724), .Q(x6_t1_w[5]) );
  DFF_X1 reg_r6_q_reg_4_ ( .D(n3636), .CK(n3724), .Q(x6_t1_w[4]) );
  DFF_X1 reg_r6_q_reg_3_ ( .D(n3652), .CK(n3724), .Q(x6_t1_w[3]) );
  DFF_X1 reg_r6_q_reg_2_ ( .D(n3668), .CK(n3724), .Q(x6_t1_w[2]) );
  DFF_X1 reg_r6_q_reg_1_ ( .D(n3684), .CK(n3724), .Q(x6_t1_w[1]) );
  DFF_X1 reg_r6_q_reg_0_ ( .D(n3700), .CK(n3724), .Q(x6_t1_w[0]) );
  DFF_X1 reg_r7_q_reg_31_ ( .D(n1000), .CK(n3724), .Q(x7_t2_w[31]) );
  DFF_X1 reg_r7_q_reg_30_ ( .D(n1016), .CK(n3724), .Q(x7_t2_w[30]) );
  DFF_X1 reg_r7_q_reg_29_ ( .D(n1032), .CK(n3724), .Q(x7_t2_w[29]) );
  DFF_X1 reg_r7_q_reg_28_ ( .D(n1048), .CK(n3724), .Q(x7_t2_w[28]) );
  DFF_X1 reg_r7_q_reg_27_ ( .D(n1064), .CK(n3724), .Q(x7_t2_w[27]) );
  DFF_X1 reg_r7_q_reg_26_ ( .D(n2639), .CK(n3724), .Q(x7_t2_w[26]) );
  DFF_X1 reg_r7_q_reg_25_ ( .D(n3301), .CK(n3724), .Q(x7_t2_w[25]) );
  DFF_X1 reg_r7_q_reg_24_ ( .D(n3317), .CK(n3724), .Q(x7_t2_w[24]) );
  DFF_X1 reg_r7_q_reg_23_ ( .D(n3333), .CK(n3724), .Q(x7_t2_w[23]) );
  DFF_X1 reg_r7_q_reg_22_ ( .D(n3349), .CK(n3724), .Q(x7_t2_w[22]) );
  DFF_X1 reg_r7_q_reg_21_ ( .D(n3365), .CK(n3724), .Q(x7_t2_w[21]) );
  DFF_X1 reg_r7_q_reg_20_ ( .D(n3381), .CK(n3724), .Q(x7_t2_w[20]) );
  DFF_X1 reg_r7_q_reg_19_ ( .D(n3397), .CK(n3724), .Q(x7_t2_w[19]) );
  DFF_X1 reg_r7_q_reg_18_ ( .D(n3413), .CK(n3724), .Q(x7_t2_w[18]) );
  DFF_X1 reg_r7_q_reg_17_ ( .D(n3429), .CK(n3724), .Q(x7_t2_w[17]) );
  DFF_X1 reg_r7_q_reg_16_ ( .D(n3445), .CK(n3724), .Q(x7_t2_w[16]) );
  DFF_X1 reg_r7_q_reg_15_ ( .D(n3461), .CK(n3724), .Q(x7_t2_w[15]) );
  DFF_X1 reg_r7_q_reg_14_ ( .D(n3477), .CK(n3724), .Q(x7_t2_w[14]) );
  DFF_X1 reg_r7_q_reg_13_ ( .D(n3493), .CK(n3724), .Q(x7_t2_w[13]) );
  DFF_X1 reg_r7_q_reg_12_ ( .D(n3509), .CK(n3724), .Q(x7_t2_w[12]) );
  DFF_X1 reg_r7_q_reg_11_ ( .D(n3525), .CK(n3724), .Q(x7_t2_w[11]) );
  DFF_X1 reg_r7_q_reg_10_ ( .D(n3541), .CK(n3724), .Q(x7_t2_w[10]) );
  DFF_X1 reg_r7_q_reg_9_ ( .D(n3557), .CK(n3724), .Q(x7_t2_w[9]) );
  DFF_X1 reg_r7_q_reg_8_ ( .D(n3573), .CK(n3724), .Q(x7_t2_w[8]) );
  DFF_X1 reg_r7_q_reg_7_ ( .D(n3589), .CK(n3724), .Q(x7_t2_w[7]) );
  DFF_X1 reg_r7_q_reg_6_ ( .D(n3605), .CK(n3724), .Q(x7_t2_w[6]) );
  DFF_X1 reg_r7_q_reg_5_ ( .D(n3621), .CK(n3724), .Q(x7_t2_w[5]) );
  DFF_X1 reg_r7_q_reg_4_ ( .D(n3637), .CK(n3724), .Q(x7_t2_w[4]) );
  DFF_X1 reg_r7_q_reg_3_ ( .D(n3653), .CK(n3724), .Q(x7_t2_w[3]) );
  DFF_X1 reg_r7_q_reg_2_ ( .D(n3669), .CK(n3724), .Q(x7_t2_w[2]) );
  DFF_X1 reg_r7_q_reg_1_ ( .D(n3685), .CK(n3724), .Q(x7_t2_w[1]) );
  DFF_X1 reg_r7_q_reg_0_ ( .D(n3701), .CK(n3724), .Q(x7_t2_w[0]) );
  DFF_X1 reg_r8_q_reg_31_ ( .D(n1001), .CK(n3724), .Q(x8_s0_w[31]) );
  DFF_X1 reg_r8_q_reg_30_ ( .D(n1017), .CK(n3724), .Q(x8_s0_w[30]) );
  DFF_X1 reg_r8_q_reg_29_ ( .D(n1033), .CK(n3724), .Q(x8_s0_w[29]) );
  DFF_X1 reg_r8_q_reg_28_ ( .D(n1049), .CK(n3724), .Q(x8_s0_w[28]) );
  DFF_X1 reg_r8_q_reg_27_ ( .D(n1065), .CK(n3724), .Q(x8_s0_w[27]) );
  DFF_X1 reg_r8_q_reg_26_ ( .D(n2640), .CK(n3724), .Q(x8_s0_w[26]) );
  DFF_X1 reg_r8_q_reg_25_ ( .D(n3302), .CK(n3724), .Q(x8_s0_w[25]) );
  DFF_X1 reg_r8_q_reg_24_ ( .D(n3318), .CK(n3724), .Q(x8_s0_w[24]) );
  DFF_X1 reg_r8_q_reg_23_ ( .D(n3334), .CK(n3724), .Q(x8_s0_w[23]) );
  DFF_X1 reg_r8_q_reg_22_ ( .D(n3350), .CK(n3724), .Q(x8_s0_w[22]) );
  DFF_X1 reg_r8_q_reg_21_ ( .D(n3366), .CK(n3724), .Q(x8_s0_w[21]) );
  DFF_X1 reg_r8_q_reg_20_ ( .D(n3382), .CK(n3724), .Q(x8_s0_w[20]) );
  DFF_X1 reg_r8_q_reg_19_ ( .D(n3398), .CK(n3724), .Q(x8_s0_w[19]) );
  DFF_X1 reg_r8_q_reg_18_ ( .D(n3414), .CK(n3724), .Q(x8_s0_w[18]) );
  DFF_X1 reg_r8_q_reg_17_ ( .D(n3430), .CK(n3724), .Q(x8_s0_w[17]) );
  DFF_X1 reg_r8_q_reg_16_ ( .D(n3446), .CK(n3724), .Q(x8_s0_w[16]) );
  DFF_X1 reg_r8_q_reg_15_ ( .D(n3462), .CK(n3724), .Q(x8_s0_w[15]) );
  DFF_X1 reg_r8_q_reg_14_ ( .D(n3478), .CK(n3724), .Q(x8_s0_w[14]) );
  DFF_X1 reg_r8_q_reg_13_ ( .D(n3494), .CK(n3724), .Q(x8_s0_w[13]) );
  DFF_X1 reg_r8_q_reg_12_ ( .D(n3510), .CK(n3724), .Q(x8_s0_w[12]) );
  DFF_X1 reg_r8_q_reg_11_ ( .D(n3526), .CK(n3724), .Q(x8_s0_w[11]) );
  DFF_X1 reg_r8_q_reg_10_ ( .D(n3542), .CK(n3724), .Q(x8_s0_w[10]) );
  DFF_X1 reg_r8_q_reg_9_ ( .D(n3558), .CK(n3724), .Q(x8_s0_w[9]) );
  DFF_X1 reg_r8_q_reg_8_ ( .D(n3574), .CK(n3724), .Q(x8_s0_w[8]) );
  DFF_X1 reg_r8_q_reg_7_ ( .D(n3590), .CK(n3724), .Q(x8_s0_w[7]) );
  DFF_X1 reg_r8_q_reg_6_ ( .D(n3606), .CK(n3724), .Q(x8_s0_w[6]) );
  DFF_X1 reg_r8_q_reg_5_ ( .D(n3622), .CK(n3724), .Q(x8_s0_w[5]) );
  DFF_X1 reg_r8_q_reg_4_ ( .D(n3638), .CK(n3724), .Q(x8_s0_w[4]) );
  DFF_X1 reg_r8_q_reg_3_ ( .D(n3654), .CK(n3724), .Q(x8_s0_w[3]) );
  DFF_X1 reg_r8_q_reg_2_ ( .D(n3670), .CK(n3724), .Q(x8_s0_w[2]) );
  DFF_X1 reg_r8_q_reg_1_ ( .D(n3686), .CK(n3724), .Q(x8_s0_w[1]) );
  DFF_X1 reg_r8_q_reg_0_ ( .D(n3702), .CK(n3724), .Q(x8_s0_w[0]) );
  DFF_X1 reg_r9_q_reg_31_ ( .D(n1002), .CK(n3724), .Q(x9_s1_w[31]) );
  DFF_X1 reg_r9_q_reg_30_ ( .D(n1018), .CK(n3724), .Q(x9_s1_w[30]) );
  DFF_X1 reg_r9_q_reg_29_ ( .D(n1034), .CK(n3724), .Q(x9_s1_w[29]) );
  DFF_X1 reg_r9_q_reg_28_ ( .D(n1050), .CK(n3724), .Q(x9_s1_w[28]) );
  DFF_X1 reg_r9_q_reg_27_ ( .D(n1066), .CK(n3724), .Q(x9_s1_w[27]) );
  DFF_X1 reg_r9_q_reg_26_ ( .D(n2641), .CK(n3724), .Q(x9_s1_w[26]) );
  DFF_X1 reg_r9_q_reg_25_ ( .D(n3303), .CK(n3724), .Q(x9_s1_w[25]) );
  DFF_X1 reg_r9_q_reg_24_ ( .D(n3319), .CK(n3724), .Q(x9_s1_w[24]) );
  DFF_X1 reg_r9_q_reg_23_ ( .D(n3335), .CK(n3724), .Q(x9_s1_w[23]) );
  DFF_X1 reg_r9_q_reg_22_ ( .D(n3351), .CK(n3724), .Q(x9_s1_w[22]) );
  DFF_X1 reg_r9_q_reg_21_ ( .D(n3367), .CK(n3724), .Q(x9_s1_w[21]) );
  DFF_X1 reg_r9_q_reg_20_ ( .D(n3383), .CK(n3724), .Q(x9_s1_w[20]) );
  DFF_X1 reg_r9_q_reg_19_ ( .D(n3399), .CK(n3724), .Q(x9_s1_w[19]) );
  DFF_X1 reg_r9_q_reg_18_ ( .D(n3415), .CK(n3724), .Q(x9_s1_w[18]) );
  DFF_X1 reg_r9_q_reg_17_ ( .D(n3431), .CK(n3724), .Q(x9_s1_w[17]) );
  DFF_X1 reg_r9_q_reg_16_ ( .D(n3447), .CK(n3724), .Q(x9_s1_w[16]) );
  DFF_X1 reg_r9_q_reg_15_ ( .D(n3463), .CK(n3724), .Q(x9_s1_w[15]) );
  DFF_X1 reg_r9_q_reg_14_ ( .D(n3479), .CK(n3724), .Q(x9_s1_w[14]) );
  DFF_X1 reg_r9_q_reg_13_ ( .D(n3495), .CK(n3724), .Q(x9_s1_w[13]) );
  DFF_X1 reg_r9_q_reg_12_ ( .D(n3511), .CK(n3724), .Q(x9_s1_w[12]) );
  DFF_X1 reg_r9_q_reg_11_ ( .D(n3527), .CK(n3724), .Q(x9_s1_w[11]) );
  DFF_X1 reg_r9_q_reg_10_ ( .D(n3543), .CK(n3724), .Q(x9_s1_w[10]) );
  DFF_X1 reg_r9_q_reg_9_ ( .D(n3559), .CK(n3724), .Q(x9_s1_w[9]) );
  DFF_X1 reg_r9_q_reg_8_ ( .D(n3575), .CK(n3724), .Q(x9_s1_w[8]) );
  DFF_X1 reg_r9_q_reg_7_ ( .D(n3591), .CK(n3724), .Q(x9_s1_w[7]) );
  DFF_X1 reg_r9_q_reg_6_ ( .D(n3607), .CK(n3724), .Q(x9_s1_w[6]) );
  DFF_X1 reg_r9_q_reg_5_ ( .D(n3623), .CK(n3724), .Q(x9_s1_w[5]) );
  DFF_X1 reg_r9_q_reg_4_ ( .D(n3639), .CK(n3724), .Q(x9_s1_w[4]) );
  DFF_X1 reg_r9_q_reg_3_ ( .D(n3655), .CK(n3724), .Q(x9_s1_w[3]) );
  DFF_X1 reg_r9_q_reg_2_ ( .D(n3671), .CK(n3724), .Q(x9_s1_w[2]) );
  DFF_X1 reg_r9_q_reg_1_ ( .D(n3687), .CK(n3724), .Q(x9_s1_w[1]) );
  DFF_X1 reg_r9_q_reg_0_ ( .D(n3703), .CK(n3724), .Q(x9_s1_w[0]) );
  DFF_X1 reg_r10_q_reg_31_ ( .D(n3098), .CK(n3724), .QN(n449) );
  DFF_X1 reg_r10_q_reg_30_ ( .D(n3097), .CK(n3724), .QN(n450) );
  DFF_X1 reg_r10_q_reg_29_ ( .D(n3096), .CK(n3724), .QN(n451) );
  DFF_X1 reg_r10_q_reg_28_ ( .D(n3095), .CK(n3724), .QN(n452) );
  DFF_X1 reg_r10_q_reg_27_ ( .D(n3094), .CK(n3724), .QN(n453) );
  DFF_X1 reg_r10_q_reg_26_ ( .D(n3093), .CK(n3724), .QN(n454) );
  DFF_X1 reg_r10_q_reg_25_ ( .D(n3092), .CK(n3724), .QN(n455) );
  DFF_X1 reg_r10_q_reg_24_ ( .D(n3091), .CK(n3724), .QN(n456) );
  DFF_X1 reg_r10_q_reg_23_ ( .D(n3090), .CK(n3724), .QN(n457) );
  DFF_X1 reg_r10_q_reg_22_ ( .D(n3089), .CK(n3724), .QN(n458) );
  DFF_X1 reg_r10_q_reg_21_ ( .D(n3088), .CK(n3724), .QN(n459) );
  DFF_X1 reg_r10_q_reg_20_ ( .D(n3087), .CK(n3724), .QN(n460) );
  DFF_X1 reg_r10_q_reg_19_ ( .D(n3086), .CK(n3724), .QN(n461) );
  DFF_X1 reg_r10_q_reg_18_ ( .D(n3085), .CK(n3724), .QN(n462) );
  DFF_X1 reg_r10_q_reg_17_ ( .D(n3084), .CK(n3724), .QN(n463) );
  DFF_X1 reg_r10_q_reg_16_ ( .D(n3083), .CK(n3724), .QN(n464) );
  DFF_X1 reg_r10_q_reg_15_ ( .D(n3082), .CK(n3724), .QN(n465) );
  DFF_X1 reg_r10_q_reg_14_ ( .D(n3081), .CK(n3724), .QN(n466) );
  DFF_X1 reg_r10_q_reg_13_ ( .D(n3080), .CK(n3724), .QN(n467) );
  DFF_X1 reg_r10_q_reg_12_ ( .D(n3079), .CK(n3724), .QN(n468) );
  DFF_X1 reg_r10_q_reg_11_ ( .D(n3078), .CK(n3724), .QN(n469) );
  DFF_X1 reg_r10_q_reg_10_ ( .D(n3077), .CK(n3724), .QN(n470) );
  DFF_X1 reg_r10_q_reg_9_ ( .D(n3076), .CK(n3724), .QN(n471) );
  DFF_X1 reg_r10_q_reg_8_ ( .D(n3075), .CK(n3724), .QN(n472) );
  DFF_X1 reg_r10_q_reg_7_ ( .D(n3074), .CK(n3724), .QN(n473) );
  DFF_X1 reg_r10_q_reg_6_ ( .D(n3073), .CK(n3724), .QN(n474) );
  DFF_X1 reg_r10_q_reg_5_ ( .D(n3072), .CK(n3724), .QN(n475) );
  DFF_X1 reg_r10_q_reg_4_ ( .D(n3071), .CK(n3724), .QN(n476) );
  DFF_X1 reg_r10_q_reg_3_ ( .D(n3070), .CK(n3724), .QN(n477) );
  DFF_X1 reg_r10_q_reg_2_ ( .D(n3069), .CK(n3724), .QN(n478) );
  DFF_X1 reg_r10_q_reg_1_ ( .D(n3068), .CK(n3724), .QN(n479) );
  DFF_X1 reg_r10_q_reg_0_ ( .D(n3067), .CK(n3724), .QN(n480) );
  DFF_X1 reg_r11_q_reg_31_ ( .D(n3066), .CK(n3724), .QN(n481) );
  DFF_X1 reg_r11_q_reg_30_ ( .D(n3065), .CK(n3724), .QN(n482) );
  DFF_X1 reg_r11_q_reg_29_ ( .D(n3064), .CK(n3724), .QN(n483) );
  DFF_X1 reg_r11_q_reg_28_ ( .D(n3063), .CK(n3724), .QN(n484) );
  DFF_X1 reg_r11_q_reg_27_ ( .D(n3062), .CK(n3724), .QN(n485) );
  DFF_X1 reg_r11_q_reg_26_ ( .D(n3061), .CK(n3724), .QN(n486) );
  DFF_X1 reg_r11_q_reg_25_ ( .D(n3060), .CK(n3724), .QN(n487) );
  DFF_X1 reg_r11_q_reg_24_ ( .D(n3059), .CK(n3724), .QN(n488) );
  DFF_X1 reg_r11_q_reg_23_ ( .D(n3058), .CK(n3724), .QN(n489) );
  DFF_X1 reg_r11_q_reg_22_ ( .D(n3057), .CK(n3724), .QN(n490) );
  DFF_X1 reg_r11_q_reg_21_ ( .D(n3056), .CK(n3724), .QN(n491) );
  DFF_X1 reg_r11_q_reg_20_ ( .D(n3055), .CK(n3724), .QN(n492) );
  DFF_X1 reg_r11_q_reg_19_ ( .D(n3054), .CK(n3724), .QN(n493) );
  DFF_X1 reg_r11_q_reg_18_ ( .D(n3053), .CK(n3724), .QN(n494) );
  DFF_X1 reg_r11_q_reg_17_ ( .D(n3052), .CK(n3724), .QN(n495) );
  DFF_X1 reg_r11_q_reg_16_ ( .D(n3051), .CK(n3724), .QN(n496) );
  DFF_X1 reg_r11_q_reg_15_ ( .D(n3050), .CK(n3724), .QN(n497) );
  DFF_X1 reg_r11_q_reg_14_ ( .D(n3049), .CK(n3724), .QN(n498) );
  DFF_X1 reg_r11_q_reg_13_ ( .D(n3048), .CK(n3724), .QN(n499) );
  DFF_X1 reg_r11_q_reg_12_ ( .D(n3047), .CK(n3724), .QN(n500) );
  DFF_X1 reg_r11_q_reg_11_ ( .D(n3046), .CK(n3724), .QN(n501) );
  DFF_X1 reg_r11_q_reg_10_ ( .D(n3045), .CK(n3724), .QN(n502) );
  DFF_X1 reg_r11_q_reg_9_ ( .D(n3044), .CK(n3724), .QN(n503) );
  DFF_X1 reg_r11_q_reg_8_ ( .D(n3043), .CK(n3724), .QN(n504) );
  DFF_X1 reg_r11_q_reg_7_ ( .D(n3042), .CK(n3724), .QN(n505) );
  DFF_X1 reg_r11_q_reg_6_ ( .D(n3041), .CK(n3724), .QN(n506) );
  DFF_X1 reg_r11_q_reg_5_ ( .D(n3040), .CK(n3724), .QN(n507) );
  DFF_X1 reg_r11_q_reg_4_ ( .D(n3039), .CK(n3724), .QN(n508) );
  DFF_X1 reg_r11_q_reg_3_ ( .D(n3038), .CK(n3724), .QN(n509) );
  DFF_X1 reg_r11_q_reg_2_ ( .D(n3037), .CK(n3724), .QN(n510) );
  DFF_X1 reg_r11_q_reg_1_ ( .D(n3036), .CK(n3724), .QN(n511) );
  DFF_X1 reg_r11_q_reg_0_ ( .D(n3035), .CK(n3724), .QN(n512) );
  DFF_X1 reg_r12_q_reg_31_ ( .D(n3034), .CK(n3724), .QN(n513) );
  DFF_X1 reg_r12_q_reg_30_ ( .D(n3033), .CK(n3724), .QN(n514) );
  DFF_X1 reg_r12_q_reg_29_ ( .D(n3032), .CK(n3724), .QN(n515) );
  DFF_X1 reg_r12_q_reg_28_ ( .D(n3031), .CK(n3724), .QN(n516) );
  DFF_X1 reg_r12_q_reg_27_ ( .D(n3030), .CK(n3724), .QN(n517) );
  DFF_X1 reg_r12_q_reg_26_ ( .D(n3029), .CK(n3724), .QN(n518) );
  DFF_X1 reg_r12_q_reg_25_ ( .D(n3028), .CK(n3724), .QN(n519) );
  DFF_X1 reg_r12_q_reg_24_ ( .D(n3027), .CK(n3724), .QN(n520) );
  DFF_X1 reg_r12_q_reg_23_ ( .D(n3026), .CK(n3724), .QN(n521) );
  DFF_X1 reg_r12_q_reg_22_ ( .D(n3025), .CK(n3724), .QN(n522) );
  DFF_X1 reg_r12_q_reg_21_ ( .D(n3024), .CK(n3724), .QN(n523) );
  DFF_X1 reg_r12_q_reg_20_ ( .D(n3023), .CK(n3724), .QN(n524) );
  DFF_X1 reg_r12_q_reg_19_ ( .D(n3022), .CK(n3724), .QN(n525) );
  DFF_X1 reg_r12_q_reg_18_ ( .D(n3021), .CK(n3724), .QN(n526) );
  DFF_X1 reg_r12_q_reg_17_ ( .D(n3020), .CK(n3724), .QN(n527) );
  DFF_X1 reg_r12_q_reg_16_ ( .D(n3019), .CK(n3724), .QN(n528) );
  DFF_X1 reg_r12_q_reg_15_ ( .D(n3018), .CK(n3724), .QN(n529) );
  DFF_X1 reg_r12_q_reg_14_ ( .D(n3017), .CK(n3724), .QN(n530) );
  DFF_X1 reg_r12_q_reg_13_ ( .D(n3016), .CK(n3724), .QN(n531) );
  DFF_X1 reg_r12_q_reg_12_ ( .D(n3015), .CK(n3724), .QN(n532) );
  DFF_X1 reg_r12_q_reg_11_ ( .D(n3014), .CK(n3724), .QN(n533) );
  DFF_X1 reg_r12_q_reg_10_ ( .D(n3013), .CK(n3724), .QN(n534) );
  DFF_X1 reg_r12_q_reg_9_ ( .D(n3012), .CK(n3724), .QN(n535) );
  DFF_X1 reg_r12_q_reg_8_ ( .D(n3011), .CK(n3724), .QN(n536) );
  DFF_X1 reg_r12_q_reg_7_ ( .D(n3010), .CK(n3724), .QN(n537) );
  DFF_X1 reg_r12_q_reg_6_ ( .D(n3009), .CK(n3724), .QN(n538) );
  DFF_X1 reg_r12_q_reg_5_ ( .D(n3008), .CK(n3724), .QN(n539) );
  DFF_X1 reg_r12_q_reg_4_ ( .D(n3007), .CK(n3724), .QN(n540) );
  DFF_X1 reg_r12_q_reg_3_ ( .D(n3006), .CK(n3724), .QN(n541) );
  DFF_X1 reg_r12_q_reg_2_ ( .D(n3005), .CK(n3724), .QN(n542) );
  DFF_X1 reg_r12_q_reg_1_ ( .D(n3004), .CK(n3724), .QN(n543) );
  DFF_X1 reg_r12_q_reg_0_ ( .D(n3003), .CK(n3724), .QN(n544) );
  DFF_X1 reg_r13_q_reg_31_ ( .D(n3002), .CK(n3724), .QN(n545) );
  DFF_X1 reg_r13_q_reg_30_ ( .D(n3001), .CK(n3724), .QN(n546) );
  DFF_X1 reg_r13_q_reg_29_ ( .D(n3000), .CK(n3724), .QN(n547) );
  DFF_X1 reg_r13_q_reg_28_ ( .D(n2999), .CK(n3724), .QN(n548) );
  DFF_X1 reg_r13_q_reg_27_ ( .D(n2998), .CK(n3724), .QN(n549) );
  DFF_X1 reg_r13_q_reg_26_ ( .D(n2997), .CK(n3724), .QN(n550) );
  DFF_X1 reg_r13_q_reg_25_ ( .D(n2996), .CK(n3724), .QN(n551) );
  DFF_X1 reg_r13_q_reg_24_ ( .D(n2995), .CK(n3724), .QN(n552) );
  DFF_X1 reg_r13_q_reg_23_ ( .D(n2994), .CK(n3724), .QN(n553) );
  DFF_X1 reg_r13_q_reg_22_ ( .D(n2993), .CK(n3724), .QN(n554) );
  DFF_X1 reg_r13_q_reg_21_ ( .D(n2992), .CK(n3724), .QN(n555) );
  DFF_X1 reg_r13_q_reg_20_ ( .D(n2991), .CK(n3724), .QN(n556) );
  DFF_X1 reg_r13_q_reg_19_ ( .D(n2990), .CK(n3724), .QN(n557) );
  DFF_X1 reg_r13_q_reg_18_ ( .D(n2989), .CK(n3724), .QN(n558) );
  DFF_X1 reg_r13_q_reg_17_ ( .D(n2988), .CK(n3724), .QN(n559) );
  DFF_X1 reg_r13_q_reg_16_ ( .D(n2987), .CK(n3724), .QN(n560) );
  DFF_X1 reg_r13_q_reg_15_ ( .D(n2986), .CK(n3724), .QN(n561) );
  DFF_X1 reg_r13_q_reg_14_ ( .D(n2985), .CK(n3724), .QN(n562) );
  DFF_X1 reg_r13_q_reg_13_ ( .D(n2984), .CK(n3724), .QN(n563) );
  DFF_X1 reg_r13_q_reg_12_ ( .D(n2983), .CK(n3724), .QN(n564) );
  DFF_X1 reg_r13_q_reg_11_ ( .D(n2982), .CK(n3724), .QN(n565) );
  DFF_X1 reg_r13_q_reg_10_ ( .D(n2981), .CK(n3724), .QN(n566) );
  DFF_X1 reg_r13_q_reg_9_ ( .D(n2980), .CK(n3724), .QN(n567) );
  DFF_X1 reg_r13_q_reg_8_ ( .D(n2979), .CK(n3724), .QN(n568) );
  DFF_X1 reg_r13_q_reg_7_ ( .D(n2978), .CK(n3724), .QN(n569) );
  DFF_X1 reg_r13_q_reg_6_ ( .D(n2977), .CK(n3724), .QN(n570) );
  DFF_X1 reg_r13_q_reg_5_ ( .D(n2976), .CK(n3724), .QN(n571) );
  DFF_X1 reg_r13_q_reg_4_ ( .D(n2975), .CK(n3724), .QN(n572) );
  DFF_X1 reg_r13_q_reg_3_ ( .D(n2974), .CK(n3724), .QN(n573) );
  DFF_X1 reg_r13_q_reg_2_ ( .D(n2973), .CK(n3724), .QN(n574) );
  DFF_X1 reg_r13_q_reg_1_ ( .D(n2972), .CK(n3724), .QN(n575) );
  DFF_X1 reg_r13_q_reg_0_ ( .D(n2971), .CK(n3724), .QN(n576) );
  DFF_X1 reg_r14_q_reg_31_ ( .D(n1003), .CK(n3724), .Q(x14_a4_w[31]) );
  DFF_X1 reg_r14_q_reg_30_ ( .D(n1019), .CK(n3724), .Q(x14_a4_w[30]) );
  DFF_X1 reg_r14_q_reg_29_ ( .D(n1035), .CK(n3724), .Q(x14_a4_w[29]) );
  DFF_X1 reg_r14_q_reg_28_ ( .D(n1051), .CK(n3724), .Q(x14_a4_w[28]) );
  DFF_X1 reg_r14_q_reg_27_ ( .D(n1067), .CK(n3724), .Q(x14_a4_w[27]) );
  DFF_X1 reg_r14_q_reg_26_ ( .D(n2643), .CK(n3724), .Q(x14_a4_w[26]) );
  DFF_X1 reg_r14_q_reg_25_ ( .D(n3304), .CK(n3724), .Q(x14_a4_w[25]) );
  DFF_X1 reg_r14_q_reg_24_ ( .D(n3320), .CK(n3724), .Q(x14_a4_w[24]) );
  DFF_X1 reg_r14_q_reg_23_ ( .D(n3336), .CK(n3724), .Q(x14_a4_w[23]) );
  DFF_X1 reg_r14_q_reg_22_ ( .D(n3352), .CK(n3724), .Q(x14_a4_w[22]) );
  DFF_X1 reg_r14_q_reg_21_ ( .D(n3368), .CK(n3724), .Q(x14_a4_w[21]) );
  DFF_X1 reg_r14_q_reg_20_ ( .D(n3384), .CK(n3724), .Q(x14_a4_w[20]) );
  DFF_X1 reg_r14_q_reg_19_ ( .D(n3400), .CK(n3724), .Q(x14_a4_w[19]) );
  DFF_X1 reg_r14_q_reg_18_ ( .D(n3416), .CK(n3724), .Q(x14_a4_w[18]) );
  DFF_X1 reg_r14_q_reg_17_ ( .D(n3432), .CK(n3724), .Q(x14_a4_w[17]) );
  DFF_X1 reg_r14_q_reg_16_ ( .D(n3448), .CK(n3724), .Q(x14_a4_w[16]) );
  DFF_X1 reg_r14_q_reg_15_ ( .D(n3464), .CK(n3724), .Q(x14_a4_w[15]) );
  DFF_X1 reg_r14_q_reg_14_ ( .D(n3480), .CK(n3724), .Q(x14_a4_w[14]) );
  DFF_X1 reg_r14_q_reg_13_ ( .D(n3496), .CK(n3724), .Q(x14_a4_w[13]) );
  DFF_X1 reg_r14_q_reg_12_ ( .D(n3512), .CK(n3724), .Q(x14_a4_w[12]) );
  DFF_X1 reg_r14_q_reg_11_ ( .D(n3528), .CK(n3724), .Q(x14_a4_w[11]) );
  DFF_X1 reg_r14_q_reg_10_ ( .D(n3544), .CK(n3724), .Q(x14_a4_w[10]) );
  DFF_X1 reg_r14_q_reg_9_ ( .D(n3560), .CK(n3724), .Q(x14_a4_w[9]) );
  DFF_X1 reg_r14_q_reg_8_ ( .D(n3576), .CK(n3724), .Q(x14_a4_w[8]) );
  DFF_X1 reg_r14_q_reg_7_ ( .D(n3592), .CK(n3724), .Q(x14_a4_w[7]) );
  DFF_X1 reg_r14_q_reg_6_ ( .D(n3608), .CK(n3724), .Q(x14_a4_w[6]) );
  DFF_X1 reg_r14_q_reg_5_ ( .D(n3624), .CK(n3724), .Q(x14_a4_w[5]) );
  DFF_X1 reg_r14_q_reg_4_ ( .D(n3640), .CK(n3724), .Q(x14_a4_w[4]) );
  DFF_X1 reg_r14_q_reg_3_ ( .D(n3656), .CK(n3724), .Q(x14_a4_w[3]) );
  DFF_X1 reg_r14_q_reg_2_ ( .D(n3672), .CK(n3724), .Q(x14_a4_w[2]) );
  DFF_X1 reg_r14_q_reg_1_ ( .D(n3688), .CK(n3724), .Q(x14_a4_w[1]) );
  DFF_X1 reg_r14_q_reg_0_ ( .D(n3704), .CK(n3724), .Q(x14_a4_w[0]) );
  DFF_X1 reg_r15_q_reg_31_ ( .D(n1004), .CK(n3724), .Q(x15_a5_w[31]) );
  DFF_X1 reg_r15_q_reg_30_ ( .D(n1020), .CK(n3724), .Q(x15_a5_w[30]) );
  DFF_X1 reg_r15_q_reg_29_ ( .D(n1036), .CK(n3724), .Q(x15_a5_w[29]) );
  DFF_X1 reg_r15_q_reg_28_ ( .D(n1052), .CK(n3724), .Q(x15_a5_w[28]) );
  DFF_X1 reg_r15_q_reg_27_ ( .D(n1068), .CK(n3724), .Q(x15_a5_w[27]) );
  DFF_X1 reg_r15_q_reg_26_ ( .D(n2777), .CK(n3724), .Q(x15_a5_w[26]) );
  DFF_X1 reg_r15_q_reg_25_ ( .D(n3305), .CK(n3724), .Q(x15_a5_w[25]) );
  DFF_X1 reg_r15_q_reg_24_ ( .D(n3321), .CK(n3724), .Q(x15_a5_w[24]) );
  DFF_X1 reg_r15_q_reg_23_ ( .D(n3337), .CK(n3724), .Q(x15_a5_w[23]) );
  DFF_X1 reg_r15_q_reg_22_ ( .D(n3353), .CK(n3724), .Q(x15_a5_w[22]) );
  DFF_X1 reg_r15_q_reg_21_ ( .D(n3369), .CK(n3724), .Q(x15_a5_w[21]) );
  DFF_X1 reg_r15_q_reg_20_ ( .D(n3385), .CK(n3724), .Q(x15_a5_w[20]) );
  DFF_X1 reg_r15_q_reg_19_ ( .D(n3401), .CK(n3724), .Q(x15_a5_w[19]) );
  DFF_X1 reg_r15_q_reg_18_ ( .D(n3417), .CK(n3724), .Q(x15_a5_w[18]) );
  DFF_X1 reg_r15_q_reg_17_ ( .D(n3433), .CK(n3724), .Q(x15_a5_w[17]) );
  DFF_X1 reg_r15_q_reg_16_ ( .D(n3449), .CK(n3724), .Q(x15_a5_w[16]) );
  DFF_X1 reg_r15_q_reg_15_ ( .D(n3465), .CK(n3724), .Q(x15_a5_w[15]) );
  DFF_X1 reg_r15_q_reg_14_ ( .D(n3481), .CK(n3724), .Q(x15_a5_w[14]) );
  DFF_X1 reg_r15_q_reg_13_ ( .D(n3497), .CK(n3724), .Q(x15_a5_w[13]) );
  DFF_X1 reg_r15_q_reg_12_ ( .D(n3513), .CK(n3724), .Q(x15_a5_w[12]) );
  DFF_X1 reg_r15_q_reg_11_ ( .D(n3529), .CK(n3724), .Q(x15_a5_w[11]) );
  DFF_X1 reg_r15_q_reg_10_ ( .D(n3545), .CK(n3724), .Q(x15_a5_w[10]) );
  DFF_X1 reg_r15_q_reg_9_ ( .D(n3561), .CK(n3724), .Q(x15_a5_w[9]) );
  DFF_X1 reg_r15_q_reg_8_ ( .D(n3577), .CK(n3724), .Q(x15_a5_w[8]) );
  DFF_X1 reg_r15_q_reg_7_ ( .D(n3593), .CK(n3724), .Q(x15_a5_w[7]) );
  DFF_X1 reg_r15_q_reg_6_ ( .D(n3609), .CK(n3724), .Q(x15_a5_w[6]) );
  DFF_X1 reg_r15_q_reg_5_ ( .D(n3625), .CK(n3724), .Q(x15_a5_w[5]) );
  DFF_X1 reg_r15_q_reg_4_ ( .D(n3641), .CK(n3724), .Q(x15_a5_w[4]) );
  DFF_X1 reg_r15_q_reg_3_ ( .D(n3657), .CK(n3724), .Q(x15_a5_w[3]) );
  DFF_X1 reg_r15_q_reg_2_ ( .D(n3673), .CK(n3724), .Q(x15_a5_w[2]) );
  DFF_X1 reg_r15_q_reg_1_ ( .D(n3689), .CK(n3724), .Q(x15_a5_w[1]) );
  DFF_X1 reg_r15_q_reg_0_ ( .D(n3705), .CK(n3724), .Q(x15_a5_w[0]) );
  DFF_X1 reg_r16_q_reg_31_ ( .D(n1005), .CK(n3724), .Q(x16_a6_w[31]) );
  DFF_X1 reg_r16_q_reg_30_ ( .D(n1021), .CK(n3724), .Q(x16_a6_w[30]) );
  DFF_X1 reg_r16_q_reg_29_ ( .D(n1037), .CK(n3724), .Q(x16_a6_w[29]) );
  DFF_X1 reg_r16_q_reg_28_ ( .D(n1053), .CK(n3724), .Q(x16_a6_w[28]) );
  DFF_X1 reg_r16_q_reg_27_ ( .D(n1069), .CK(n3724), .Q(x16_a6_w[27]) );
  DFF_X1 reg_r16_q_reg_26_ ( .D(n2778), .CK(n3724), .Q(x16_a6_w[26]) );
  DFF_X1 reg_r16_q_reg_25_ ( .D(n3306), .CK(n3724), .Q(x16_a6_w[25]) );
  DFF_X1 reg_r16_q_reg_24_ ( .D(n3322), .CK(n3724), .Q(x16_a6_w[24]) );
  DFF_X1 reg_r16_q_reg_23_ ( .D(n3338), .CK(n3724), .Q(x16_a6_w[23]) );
  DFF_X1 reg_r16_q_reg_22_ ( .D(n3354), .CK(n3724), .Q(x16_a6_w[22]) );
  DFF_X1 reg_r16_q_reg_21_ ( .D(n3370), .CK(n3724), .Q(x16_a6_w[21]) );
  DFF_X1 reg_r16_q_reg_20_ ( .D(n3386), .CK(n3724), .Q(x16_a6_w[20]) );
  DFF_X1 reg_r16_q_reg_19_ ( .D(n3402), .CK(n3724), .Q(x16_a6_w[19]) );
  DFF_X1 reg_r16_q_reg_18_ ( .D(n3418), .CK(n3724), .Q(x16_a6_w[18]) );
  DFF_X1 reg_r16_q_reg_17_ ( .D(n3434), .CK(n3724), .Q(x16_a6_w[17]) );
  DFF_X1 reg_r16_q_reg_16_ ( .D(n3450), .CK(n3724), .Q(x16_a6_w[16]) );
  DFF_X1 reg_r16_q_reg_15_ ( .D(n3466), .CK(n3724), .Q(x16_a6_w[15]) );
  DFF_X1 reg_r16_q_reg_14_ ( .D(n3482), .CK(n3724), .Q(x16_a6_w[14]) );
  DFF_X1 reg_r16_q_reg_13_ ( .D(n3498), .CK(n3724), .Q(x16_a6_w[13]) );
  DFF_X1 reg_r16_q_reg_12_ ( .D(n3514), .CK(n3724), .Q(x16_a6_w[12]) );
  DFF_X1 reg_r16_q_reg_11_ ( .D(n3530), .CK(n3724), .Q(x16_a6_w[11]) );
  DFF_X1 reg_r16_q_reg_10_ ( .D(n3546), .CK(n3724), .Q(x16_a6_w[10]) );
  DFF_X1 reg_r16_q_reg_9_ ( .D(n3562), .CK(n3724), .Q(x16_a6_w[9]) );
  DFF_X1 reg_r16_q_reg_8_ ( .D(n3578), .CK(n3724), .Q(x16_a6_w[8]) );
  DFF_X1 reg_r16_q_reg_7_ ( .D(n3594), .CK(n3724), .Q(x16_a6_w[7]) );
  DFF_X1 reg_r16_q_reg_6_ ( .D(n3610), .CK(n3724), .Q(x16_a6_w[6]) );
  DFF_X1 reg_r16_q_reg_5_ ( .D(n3626), .CK(n3724), .Q(x16_a6_w[5]) );
  DFF_X1 reg_r16_q_reg_4_ ( .D(n3642), .CK(n3724), .Q(x16_a6_w[4]) );
  DFF_X1 reg_r16_q_reg_3_ ( .D(n3658), .CK(n3724), .Q(x16_a6_w[3]) );
  DFF_X1 reg_r16_q_reg_2_ ( .D(n3674), .CK(n3724), .Q(x16_a6_w[2]) );
  DFF_X1 reg_r16_q_reg_1_ ( .D(n3690), .CK(n3724), .Q(x16_a6_w[1]) );
  DFF_X1 reg_r16_q_reg_0_ ( .D(n3706), .CK(n3724), .Q(x16_a6_w[0]) );
  DFF_X1 reg_r17_q_reg_31_ ( .D(n1006), .CK(n3724), .Q(x17_a7_w[31]) );
  DFF_X1 reg_r17_q_reg_30_ ( .D(n1022), .CK(n3724), .Q(x17_a7_w[30]) );
  DFF_X1 reg_r17_q_reg_29_ ( .D(n1038), .CK(n3724), .Q(x17_a7_w[29]) );
  DFF_X1 reg_r17_q_reg_28_ ( .D(n1054), .CK(n3724), .Q(x17_a7_w[28]) );
  DFF_X1 reg_r17_q_reg_27_ ( .D(n2285), .CK(n3724), .Q(x17_a7_w[27]) );
  DFF_X1 reg_r17_q_reg_26_ ( .D(n3291), .CK(n3724), .Q(x17_a7_w[26]) );
  DFF_X1 reg_r17_q_reg_25_ ( .D(n3307), .CK(n3724), .Q(x17_a7_w[25]) );
  DFF_X1 reg_r17_q_reg_24_ ( .D(n3323), .CK(n3724), .Q(x17_a7_w[24]) );
  DFF_X1 reg_r17_q_reg_23_ ( .D(n3339), .CK(n3724), .Q(x17_a7_w[23]) );
  DFF_X1 reg_r17_q_reg_22_ ( .D(n3355), .CK(n3724), .Q(x17_a7_w[22]) );
  DFF_X1 reg_r17_q_reg_21_ ( .D(n3371), .CK(n3724), .Q(x17_a7_w[21]) );
  DFF_X1 reg_r17_q_reg_20_ ( .D(n3387), .CK(n3724), .Q(x17_a7_w[20]) );
  DFF_X1 reg_r17_q_reg_19_ ( .D(n3403), .CK(n3724), .Q(x17_a7_w[19]) );
  DFF_X1 reg_r17_q_reg_18_ ( .D(n3419), .CK(n3724), .Q(x17_a7_w[18]) );
  DFF_X1 reg_r17_q_reg_17_ ( .D(n3435), .CK(n3724), .Q(x17_a7_w[17]) );
  DFF_X1 reg_r17_q_reg_16_ ( .D(n3451), .CK(n3724), .Q(x17_a7_w[16]) );
  DFF_X1 reg_r17_q_reg_15_ ( .D(n3467), .CK(n3724), .Q(x17_a7_w[15]) );
  DFF_X1 reg_r17_q_reg_14_ ( .D(n3483), .CK(n3724), .Q(x17_a7_w[14]) );
  DFF_X1 reg_r17_q_reg_13_ ( .D(n3499), .CK(n3724), .Q(x17_a7_w[13]) );
  DFF_X1 reg_r17_q_reg_12_ ( .D(n3515), .CK(n3724), .Q(x17_a7_w[12]) );
  DFF_X1 reg_r17_q_reg_11_ ( .D(n3531), .CK(n3724), .Q(x17_a7_w[11]) );
  DFF_X1 reg_r17_q_reg_10_ ( .D(n3547), .CK(n3724), .Q(x17_a7_w[10]) );
  DFF_X1 reg_r17_q_reg_9_ ( .D(n3563), .CK(n3724), .Q(x17_a7_w[9]) );
  DFF_X1 reg_r17_q_reg_8_ ( .D(n3579), .CK(n3724), .Q(x17_a7_w[8]) );
  DFF_X1 reg_r17_q_reg_7_ ( .D(n3595), .CK(n3724), .Q(x17_a7_w[7]) );
  DFF_X1 reg_r17_q_reg_6_ ( .D(n3611), .CK(n3724), .Q(x17_a7_w[6]) );
  DFF_X1 reg_r17_q_reg_5_ ( .D(n3627), .CK(n3724), .Q(x17_a7_w[5]) );
  DFF_X1 reg_r17_q_reg_4_ ( .D(n3643), .CK(n3724), .Q(x17_a7_w[4]) );
  DFF_X1 reg_r17_q_reg_3_ ( .D(n3659), .CK(n3724), .Q(x17_a7_w[3]) );
  DFF_X1 reg_r17_q_reg_2_ ( .D(n3675), .CK(n3724), .Q(x17_a7_w[2]) );
  DFF_X1 reg_r17_q_reg_1_ ( .D(n3691), .CK(n3724), .Q(x17_a7_w[1]) );
  DFF_X1 reg_r17_q_reg_0_ ( .D(n3707), .CK(n3724), .Q(x17_a7_w[0]) );
  DFF_X1 reg_r18_q_reg_31_ ( .D(n2970), .CK(n3724), .QN(n705) );
  DFF_X1 reg_r18_q_reg_30_ ( .D(n2969), .CK(n3724), .QN(n706) );
  DFF_X1 reg_r18_q_reg_29_ ( .D(n2968), .CK(n3724), .QN(n707) );
  DFF_X1 reg_r18_q_reg_28_ ( .D(n2967), .CK(n3724), .QN(n708) );
  DFF_X1 reg_r18_q_reg_27_ ( .D(n2966), .CK(n3724), .QN(n709) );
  DFF_X1 reg_r18_q_reg_26_ ( .D(n2965), .CK(n3724), .QN(n710) );
  DFF_X1 reg_r18_q_reg_25_ ( .D(n2964), .CK(n3724), .QN(n711) );
  DFF_X1 reg_r18_q_reg_24_ ( .D(n2963), .CK(n3724), .QN(n712) );
  DFF_X1 reg_r18_q_reg_23_ ( .D(n2962), .CK(n3724), .QN(n713) );
  DFF_X1 reg_r18_q_reg_22_ ( .D(n2961), .CK(n3724), .QN(n714) );
  DFF_X1 reg_r18_q_reg_21_ ( .D(n2960), .CK(n3724), .QN(n715) );
  DFF_X1 reg_r18_q_reg_20_ ( .D(n2959), .CK(n3724), .QN(n716) );
  DFF_X1 reg_r18_q_reg_19_ ( .D(n2958), .CK(n3724), .QN(n717) );
  DFF_X1 reg_r18_q_reg_18_ ( .D(n2957), .CK(n3724), .QN(n718) );
  DFF_X1 reg_r18_q_reg_17_ ( .D(n2956), .CK(n3724), .QN(n719) );
  DFF_X1 reg_r18_q_reg_16_ ( .D(n2955), .CK(n3724), .QN(n720) );
  DFF_X1 reg_r18_q_reg_15_ ( .D(n2954), .CK(n3724), .QN(n721) );
  DFF_X1 reg_r18_q_reg_14_ ( .D(n2953), .CK(n3724), .QN(n722) );
  DFF_X1 reg_r18_q_reg_13_ ( .D(n2952), .CK(n3724), .QN(n723) );
  DFF_X1 reg_r18_q_reg_12_ ( .D(n2951), .CK(n3724), .QN(n724) );
  DFF_X1 reg_r18_q_reg_11_ ( .D(n2950), .CK(n3724), .QN(n725) );
  DFF_X1 reg_r18_q_reg_10_ ( .D(n2949), .CK(n3724), .QN(n726) );
  DFF_X1 reg_r18_q_reg_9_ ( .D(n2948), .CK(n3724), .QN(n727) );
  DFF_X1 reg_r18_q_reg_8_ ( .D(n2947), .CK(n3724), .QN(n728) );
  DFF_X1 reg_r18_q_reg_7_ ( .D(n2946), .CK(n3724), .QN(n729) );
  DFF_X1 reg_r18_q_reg_6_ ( .D(n2945), .CK(n3724), .QN(n730) );
  DFF_X1 reg_r18_q_reg_5_ ( .D(n2944), .CK(n3724), .QN(n731) );
  DFF_X1 reg_r18_q_reg_4_ ( .D(n2943), .CK(n3724), .QN(n732) );
  DFF_X1 reg_r18_q_reg_3_ ( .D(n2942), .CK(n3724), .QN(n733) );
  DFF_X1 reg_r18_q_reg_2_ ( .D(n2941), .CK(n3724), .QN(n734) );
  DFF_X1 reg_r18_q_reg_1_ ( .D(n2940), .CK(n3724), .QN(n735) );
  DFF_X1 reg_r18_q_reg_0_ ( .D(n2939), .CK(n3724), .QN(n736) );
  DFF_X1 reg_r19_q_reg_31_ ( .D(n2938), .CK(n3724), .QN(n737) );
  DFF_X1 reg_r19_q_reg_30_ ( .D(n2937), .CK(n3724), .QN(n738) );
  DFF_X1 reg_r19_q_reg_29_ ( .D(n2936), .CK(n3724), .QN(n739) );
  DFF_X1 reg_r19_q_reg_28_ ( .D(n2935), .CK(n3724), .QN(n740) );
  DFF_X1 reg_r19_q_reg_27_ ( .D(n2934), .CK(n3724), .QN(n741) );
  DFF_X1 reg_r19_q_reg_26_ ( .D(n2933), .CK(n3724), .QN(n742) );
  DFF_X1 reg_r19_q_reg_25_ ( .D(n2932), .CK(n3724), .QN(n743) );
  DFF_X1 reg_r19_q_reg_24_ ( .D(n2931), .CK(n3724), .QN(n744) );
  DFF_X1 reg_r19_q_reg_23_ ( .D(n2930), .CK(n3724), .QN(n745) );
  DFF_X1 reg_r19_q_reg_22_ ( .D(n2929), .CK(n3724), .QN(n746) );
  DFF_X1 reg_r19_q_reg_21_ ( .D(n2928), .CK(n3724), .QN(n747) );
  DFF_X1 reg_r19_q_reg_20_ ( .D(n2927), .CK(n3724), .QN(n748) );
  DFF_X1 reg_r19_q_reg_19_ ( .D(n2926), .CK(n3724), .QN(n749) );
  DFF_X1 reg_r19_q_reg_18_ ( .D(n2925), .CK(n3724), .QN(n750) );
  DFF_X1 reg_r19_q_reg_17_ ( .D(n2924), .CK(n3724), .QN(n751) );
  DFF_X1 reg_r19_q_reg_16_ ( .D(n2923), .CK(n3724), .QN(n752) );
  DFF_X1 reg_r19_q_reg_15_ ( .D(n2922), .CK(n3724), .QN(n753) );
  DFF_X1 reg_r19_q_reg_14_ ( .D(n2921), .CK(n3724), .QN(n754) );
  DFF_X1 reg_r19_q_reg_13_ ( .D(n2920), .CK(n3724), .QN(n755) );
  DFF_X1 reg_r19_q_reg_12_ ( .D(n2919), .CK(n3724), .QN(n756) );
  DFF_X1 reg_r19_q_reg_11_ ( .D(n2918), .CK(n3724), .QN(n757) );
  DFF_X1 reg_r19_q_reg_10_ ( .D(n2917), .CK(n3724), .QN(n758) );
  DFF_X1 reg_r19_q_reg_9_ ( .D(n2916), .CK(n3724), .QN(n759) );
  DFF_X1 reg_r19_q_reg_8_ ( .D(n2915), .CK(n3724), .QN(n760) );
  DFF_X1 reg_r19_q_reg_7_ ( .D(n2914), .CK(n3724), .QN(n761) );
  DFF_X1 reg_r19_q_reg_6_ ( .D(n2913), .CK(n3724), .QN(n762) );
  DFF_X1 reg_r19_q_reg_5_ ( .D(n2912), .CK(n3724), .QN(n763) );
  DFF_X1 reg_r19_q_reg_4_ ( .D(n2911), .CK(n3724), .QN(n764) );
  DFF_X1 reg_r19_q_reg_3_ ( .D(n2910), .CK(n3724), .QN(n765) );
  DFF_X1 reg_r19_q_reg_2_ ( .D(n2909), .CK(n3724), .QN(n766) );
  DFF_X1 reg_r19_q_reg_1_ ( .D(n2908), .CK(n3724), .QN(n767) );
  DFF_X1 reg_r19_q_reg_0_ ( .D(n2907), .CK(n3724), .QN(n768) );
  DFF_X1 reg_r20_q_reg_31_ ( .D(n2906), .CK(n3724), .QN(n769) );
  DFF_X1 reg_r20_q_reg_30_ ( .D(n2905), .CK(n3724), .QN(n770) );
  DFF_X1 reg_r20_q_reg_29_ ( .D(n2904), .CK(n3724), .QN(n771) );
  DFF_X1 reg_r20_q_reg_28_ ( .D(n2903), .CK(n3724), .QN(n772) );
  DFF_X1 reg_r20_q_reg_27_ ( .D(n2902), .CK(n3724), .QN(n773) );
  DFF_X1 reg_r20_q_reg_26_ ( .D(n2901), .CK(n3724), .QN(n774) );
  DFF_X1 reg_r20_q_reg_25_ ( .D(n2900), .CK(n3724), .QN(n775) );
  DFF_X1 reg_r20_q_reg_24_ ( .D(n2899), .CK(n3724), .QN(n776) );
  DFF_X1 reg_r20_q_reg_23_ ( .D(n2898), .CK(n3724), .QN(n777) );
  DFF_X1 reg_r20_q_reg_22_ ( .D(n2897), .CK(n3724), .QN(n778) );
  DFF_X1 reg_r20_q_reg_21_ ( .D(n2896), .CK(n3724), .QN(n779) );
  DFF_X1 reg_r20_q_reg_20_ ( .D(n2895), .CK(n3724), .QN(n780) );
  DFF_X1 reg_r20_q_reg_19_ ( .D(n2894), .CK(n3724), .QN(n781) );
  DFF_X1 reg_r20_q_reg_18_ ( .D(n2893), .CK(n3724), .QN(n782) );
  DFF_X1 reg_r20_q_reg_17_ ( .D(n2892), .CK(n3724), .QN(n783) );
  DFF_X1 reg_r20_q_reg_16_ ( .D(n2891), .CK(n3724), .QN(n784) );
  DFF_X1 reg_r20_q_reg_15_ ( .D(n2890), .CK(n3724), .QN(n785) );
  DFF_X1 reg_r20_q_reg_14_ ( .D(n2889), .CK(n3724), .QN(n786) );
  DFF_X1 reg_r20_q_reg_13_ ( .D(n2888), .CK(n3724), .QN(n787) );
  DFF_X1 reg_r20_q_reg_12_ ( .D(n2887), .CK(n3724), .QN(n788) );
  DFF_X1 reg_r20_q_reg_11_ ( .D(n2886), .CK(n3724), .QN(n789) );
  DFF_X1 reg_r20_q_reg_10_ ( .D(n2885), .CK(n3724), .QN(n790) );
  DFF_X1 reg_r20_q_reg_9_ ( .D(n2884), .CK(n3724), .QN(n791) );
  DFF_X1 reg_r20_q_reg_8_ ( .D(n2883), .CK(n3724), .QN(n792) );
  DFF_X1 reg_r20_q_reg_7_ ( .D(n2882), .CK(n3724), .QN(n793) );
  DFF_X1 reg_r20_q_reg_6_ ( .D(n2881), .CK(n3724), .QN(n794) );
  DFF_X1 reg_r20_q_reg_5_ ( .D(n2880), .CK(n3724), .QN(n795) );
  DFF_X1 reg_r20_q_reg_4_ ( .D(n2879), .CK(n3724), .QN(n796) );
  DFF_X1 reg_r20_q_reg_3_ ( .D(n2878), .CK(n3724), .QN(n797) );
  DFF_X1 reg_r20_q_reg_2_ ( .D(n2877), .CK(n3724), .QN(n798) );
  DFF_X1 reg_r20_q_reg_1_ ( .D(n2876), .CK(n3724), .QN(n799) );
  DFF_X1 reg_r20_q_reg_0_ ( .D(n2875), .CK(n3724), .QN(n800) );
  DFF_X1 reg_r21_q_reg_31_ ( .D(n2874), .CK(n3724), .QN(n801) );
  DFF_X1 reg_r21_q_reg_30_ ( .D(n2873), .CK(n3724), .QN(n802) );
  DFF_X1 reg_r21_q_reg_29_ ( .D(n2872), .CK(n3724), .QN(n803) );
  DFF_X1 reg_r21_q_reg_28_ ( .D(n2871), .CK(n3724), .QN(n804) );
  DFF_X1 reg_r21_q_reg_27_ ( .D(n2870), .CK(n3724), .QN(n805) );
  DFF_X1 reg_r21_q_reg_26_ ( .D(n2869), .CK(n3724), .QN(n806) );
  DFF_X1 reg_r21_q_reg_25_ ( .D(n2868), .CK(n3724), .QN(n807) );
  DFF_X1 reg_r21_q_reg_24_ ( .D(n2867), .CK(n3724), .QN(n808) );
  DFF_X1 reg_r21_q_reg_23_ ( .D(n2866), .CK(n3724), .QN(n809) );
  DFF_X1 reg_r21_q_reg_22_ ( .D(n2865), .CK(n3724), .QN(n810) );
  DFF_X1 reg_r21_q_reg_21_ ( .D(n2864), .CK(n3724), .QN(n811) );
  DFF_X1 reg_r21_q_reg_20_ ( .D(n2863), .CK(n3724), .QN(n812) );
  DFF_X1 reg_r21_q_reg_19_ ( .D(n2862), .CK(n3724), .QN(n813) );
  DFF_X1 reg_r21_q_reg_18_ ( .D(n2861), .CK(n3724), .QN(n814) );
  DFF_X1 reg_r21_q_reg_17_ ( .D(n2860), .CK(n3724), .QN(n815) );
  DFF_X1 reg_r21_q_reg_16_ ( .D(n2859), .CK(n3724), .QN(n816) );
  DFF_X1 reg_r21_q_reg_15_ ( .D(n2858), .CK(n3724), .QN(n817) );
  DFF_X1 reg_r21_q_reg_14_ ( .D(n2857), .CK(n3724), .QN(n818) );
  DFF_X1 reg_r21_q_reg_13_ ( .D(n2856), .CK(n3724), .QN(n819) );
  DFF_X1 reg_r21_q_reg_12_ ( .D(n2855), .CK(n3724), .QN(n820) );
  DFF_X1 reg_r21_q_reg_11_ ( .D(n2854), .CK(n3724), .QN(n821) );
  DFF_X1 reg_r21_q_reg_10_ ( .D(n2853), .CK(n3724), .QN(n822) );
  DFF_X1 reg_r21_q_reg_9_ ( .D(n2852), .CK(n3724), .QN(n823) );
  DFF_X1 reg_r21_q_reg_8_ ( .D(n2851), .CK(n3724), .QN(n824) );
  DFF_X1 reg_r21_q_reg_7_ ( .D(n2850), .CK(n3724), .QN(n825) );
  DFF_X1 reg_r21_q_reg_6_ ( .D(n2849), .CK(n3724), .QN(n826) );
  DFF_X1 reg_r21_q_reg_5_ ( .D(n2848), .CK(n3724), .QN(n827) );
  DFF_X1 reg_r21_q_reg_4_ ( .D(n2847), .CK(n3724), .QN(n828) );
  DFF_X1 reg_r21_q_reg_3_ ( .D(n2846), .CK(n3724), .QN(n829) );
  DFF_X1 reg_r21_q_reg_2_ ( .D(n2845), .CK(n3724), .QN(n830) );
  DFF_X1 reg_r21_q_reg_1_ ( .D(n2844), .CK(n3724), .QN(n831) );
  DFF_X1 reg_r21_q_reg_0_ ( .D(n2843), .CK(n3724), .QN(n832) );
  DFF_X1 reg_r22_q_reg_31_ ( .D(n1007), .CK(n3724), .Q(x22_s6_w[31]) );
  DFF_X1 reg_r22_q_reg_30_ ( .D(n1023), .CK(n3724), .Q(x22_s6_w[30]) );
  DFF_X1 reg_r22_q_reg_29_ ( .D(n1039), .CK(n3724), .Q(x22_s6_w[29]) );
  DFF_X1 reg_r22_q_reg_28_ ( .D(n1055), .CK(n3724), .Q(x22_s6_w[28]) );
  DFF_X1 reg_r22_q_reg_27_ ( .D(n2287), .CK(n3724), .Q(x22_s6_w[27]) );
  DFF_X1 reg_r22_q_reg_26_ ( .D(n3292), .CK(n3724), .Q(x22_s6_w[26]) );
  DFF_X1 reg_r22_q_reg_25_ ( .D(n3308), .CK(n3724), .Q(x22_s6_w[25]) );
  DFF_X1 reg_r22_q_reg_24_ ( .D(n3324), .CK(n3724), .Q(x22_s6_w[24]) );
  DFF_X1 reg_r22_q_reg_23_ ( .D(n3340), .CK(n3724), .Q(x22_s6_w[23]) );
  DFF_X1 reg_r22_q_reg_22_ ( .D(n3356), .CK(n3724), .Q(x22_s6_w[22]) );
  DFF_X1 reg_r22_q_reg_21_ ( .D(n3372), .CK(n3724), .Q(x22_s6_w[21]) );
  DFF_X1 reg_r22_q_reg_20_ ( .D(n3388), .CK(n3724), .Q(x22_s6_w[20]) );
  DFF_X1 reg_r22_q_reg_19_ ( .D(n3404), .CK(n3724), .Q(x22_s6_w[19]) );
  DFF_X1 reg_r22_q_reg_18_ ( .D(n3420), .CK(n3724), .Q(x22_s6_w[18]) );
  DFF_X1 reg_r22_q_reg_17_ ( .D(n3436), .CK(n3724), .Q(x22_s6_w[17]) );
  DFF_X1 reg_r22_q_reg_16_ ( .D(n3452), .CK(n3724), .Q(x22_s6_w[16]) );
  DFF_X1 reg_r22_q_reg_15_ ( .D(n3468), .CK(n3724), .Q(x22_s6_w[15]) );
  DFF_X1 reg_r22_q_reg_14_ ( .D(n3484), .CK(n3724), .Q(x22_s6_w[14]) );
  DFF_X1 reg_r22_q_reg_13_ ( .D(n3500), .CK(n3724), .Q(x22_s6_w[13]) );
  DFF_X1 reg_r22_q_reg_12_ ( .D(n3516), .CK(n3724), .Q(x22_s6_w[12]) );
  DFF_X1 reg_r22_q_reg_11_ ( .D(n3532), .CK(n3724), .Q(x22_s6_w[11]) );
  DFF_X1 reg_r22_q_reg_10_ ( .D(n3548), .CK(n3724), .Q(x22_s6_w[10]) );
  DFF_X1 reg_r22_q_reg_9_ ( .D(n3564), .CK(n3724), .Q(x22_s6_w[9]) );
  DFF_X1 reg_r22_q_reg_8_ ( .D(n3580), .CK(n3724), .Q(x22_s6_w[8]) );
  DFF_X1 reg_r22_q_reg_7_ ( .D(n3596), .CK(n3724), .Q(x22_s6_w[7]) );
  DFF_X1 reg_r22_q_reg_6_ ( .D(n3612), .CK(n3724), .Q(x22_s6_w[6]) );
  DFF_X1 reg_r22_q_reg_5_ ( .D(n3628), .CK(n3724), .Q(x22_s6_w[5]) );
  DFF_X1 reg_r22_q_reg_4_ ( .D(n3644), .CK(n3724), .Q(x22_s6_w[4]) );
  DFF_X1 reg_r22_q_reg_3_ ( .D(n3660), .CK(n3724), .Q(x22_s6_w[3]) );
  DFF_X1 reg_r22_q_reg_2_ ( .D(n3676), .CK(n3724), .Q(x22_s6_w[2]) );
  DFF_X1 reg_r22_q_reg_1_ ( .D(n3692), .CK(n3724), .Q(x22_s6_w[1]) );
  DFF_X1 reg_r22_q_reg_0_ ( .D(n3708), .CK(n3724), .Q(x22_s6_w[0]) );
  DFF_X1 reg_r23_q_reg_31_ ( .D(n1008), .CK(n3724), .Q(x23_s7_w[31]) );
  DFF_X1 reg_r23_q_reg_30_ ( .D(n1024), .CK(n3724), .Q(x23_s7_w[30]) );
  DFF_X1 reg_r23_q_reg_29_ ( .D(n1040), .CK(n3724), .Q(x23_s7_w[29]) );
  DFF_X1 reg_r23_q_reg_28_ ( .D(n1056), .CK(n3724), .Q(x23_s7_w[28]) );
  DFF_X1 reg_r23_q_reg_27_ ( .D(n2357), .CK(n3724), .Q(x23_s7_w[27]) );
  DFF_X1 reg_r23_q_reg_26_ ( .D(n3293), .CK(n3724), .Q(x23_s7_w[26]) );
  DFF_X1 reg_r23_q_reg_25_ ( .D(n3309), .CK(n3724), .Q(x23_s7_w[25]) );
  DFF_X1 reg_r23_q_reg_24_ ( .D(n3325), .CK(n3724), .Q(x23_s7_w[24]) );
  DFF_X1 reg_r23_q_reg_23_ ( .D(n3341), .CK(n3724), .Q(x23_s7_w[23]) );
  DFF_X1 reg_r23_q_reg_22_ ( .D(n3357), .CK(n3724), .Q(x23_s7_w[22]) );
  DFF_X1 reg_r23_q_reg_21_ ( .D(n3373), .CK(n3724), .Q(x23_s7_w[21]) );
  DFF_X1 reg_r23_q_reg_20_ ( .D(n3389), .CK(n3724), .Q(x23_s7_w[20]) );
  DFF_X1 reg_r23_q_reg_19_ ( .D(n3405), .CK(n3724), .Q(x23_s7_w[19]) );
  DFF_X1 reg_r23_q_reg_18_ ( .D(n3421), .CK(n3724), .Q(x23_s7_w[18]) );
  DFF_X1 reg_r23_q_reg_17_ ( .D(n3437), .CK(n3724), .Q(x23_s7_w[17]) );
  DFF_X1 reg_r23_q_reg_16_ ( .D(n3453), .CK(n3724), .Q(x23_s7_w[16]) );
  DFF_X1 reg_r23_q_reg_15_ ( .D(n3469), .CK(n3724), .Q(x23_s7_w[15]) );
  DFF_X1 reg_r23_q_reg_14_ ( .D(n3485), .CK(n3724), .Q(x23_s7_w[14]) );
  DFF_X1 reg_r23_q_reg_13_ ( .D(n3501), .CK(n3724), .Q(x23_s7_w[13]) );
  DFF_X1 reg_r23_q_reg_12_ ( .D(n3517), .CK(n3724), .Q(x23_s7_w[12]) );
  DFF_X1 reg_r23_q_reg_11_ ( .D(n3533), .CK(n3724), .Q(x23_s7_w[11]) );
  DFF_X1 reg_r23_q_reg_10_ ( .D(n3549), .CK(n3724), .Q(x23_s7_w[10]) );
  DFF_X1 reg_r23_q_reg_9_ ( .D(n3565), .CK(n3724), .Q(x23_s7_w[9]) );
  DFF_X1 reg_r23_q_reg_8_ ( .D(n3581), .CK(n3724), .Q(x23_s7_w[8]) );
  DFF_X1 reg_r23_q_reg_7_ ( .D(n3597), .CK(n3724), .Q(x23_s7_w[7]) );
  DFF_X1 reg_r23_q_reg_6_ ( .D(n3613), .CK(n3724), .Q(x23_s7_w[6]) );
  DFF_X1 reg_r23_q_reg_5_ ( .D(n3629), .CK(n3724), .Q(x23_s7_w[5]) );
  DFF_X1 reg_r23_q_reg_4_ ( .D(n3645), .CK(n3724), .Q(x23_s7_w[4]) );
  DFF_X1 reg_r23_q_reg_3_ ( .D(n3661), .CK(n3724), .Q(x23_s7_w[3]) );
  DFF_X1 reg_r23_q_reg_2_ ( .D(n3677), .CK(n3724), .Q(x23_s7_w[2]) );
  DFF_X1 reg_r23_q_reg_1_ ( .D(n3693), .CK(n3724), .Q(x23_s7_w[1]) );
  DFF_X1 reg_r23_q_reg_0_ ( .D(n3709), .CK(n3724), .Q(x23_s7_w[0]) );
  DFF_X1 reg_r24_q_reg_31_ ( .D(n2842), .CK(n3724), .QN(n897) );
  DFF_X1 reg_r24_q_reg_30_ ( .D(n2841), .CK(n3724), .QN(n898) );
  DFF_X1 reg_r24_q_reg_29_ ( .D(n2840), .CK(n3724), .QN(n899) );
  DFF_X1 reg_r24_q_reg_28_ ( .D(n2839), .CK(n3724), .QN(n900) );
  DFF_X1 reg_r24_q_reg_27_ ( .D(n2838), .CK(n3724), .QN(n901) );
  DFF_X1 reg_r24_q_reg_26_ ( .D(n2837), .CK(n3724), .QN(n902) );
  DFF_X1 reg_r24_q_reg_25_ ( .D(n2836), .CK(n3724), .QN(n903) );
  DFF_X1 reg_r24_q_reg_24_ ( .D(n2835), .CK(n3724), .QN(n904) );
  DFF_X1 reg_r24_q_reg_23_ ( .D(n2834), .CK(n3724), .QN(n905) );
  DFF_X1 reg_r24_q_reg_22_ ( .D(n2833), .CK(n3724), .QN(n906) );
  DFF_X1 reg_r24_q_reg_21_ ( .D(n2832), .CK(n3724), .QN(n907) );
  DFF_X1 reg_r24_q_reg_20_ ( .D(n2831), .CK(n3724), .QN(n908) );
  DFF_X1 reg_r24_q_reg_19_ ( .D(n2830), .CK(n3724), .QN(n909) );
  DFF_X1 reg_r24_q_reg_18_ ( .D(n2829), .CK(n3724), .QN(n910) );
  DFF_X1 reg_r24_q_reg_17_ ( .D(n2828), .CK(n3724), .QN(n911) );
  DFF_X1 reg_r24_q_reg_16_ ( .D(n2827), .CK(n3724), .QN(n912) );
  DFF_X1 reg_r24_q_reg_15_ ( .D(n2826), .CK(n3724), .QN(n913) );
  DFF_X1 reg_r24_q_reg_14_ ( .D(n2825), .CK(n3724), .QN(n914) );
  DFF_X1 reg_r24_q_reg_13_ ( .D(n2824), .CK(n3724), .QN(n915) );
  DFF_X1 reg_r24_q_reg_12_ ( .D(n2823), .CK(n3724), .QN(n916) );
  DFF_X1 reg_r24_q_reg_11_ ( .D(n2822), .CK(n3724), .QN(n917) );
  DFF_X1 reg_r24_q_reg_10_ ( .D(n2821), .CK(n3724), .QN(n918) );
  DFF_X1 reg_r24_q_reg_9_ ( .D(n2820), .CK(n3724), .QN(n919) );
  DFF_X1 reg_r24_q_reg_8_ ( .D(n2819), .CK(n3724), .QN(n920) );
  DFF_X1 reg_r24_q_reg_7_ ( .D(n2818), .CK(n3724), .QN(n921) );
  DFF_X1 reg_r24_q_reg_6_ ( .D(n2817), .CK(n3724), .QN(n922) );
  DFF_X1 reg_r24_q_reg_5_ ( .D(n2816), .CK(n3724), .QN(n923) );
  DFF_X1 reg_r24_q_reg_4_ ( .D(n2815), .CK(n3724), .QN(n924) );
  DFF_X1 reg_r24_q_reg_3_ ( .D(n2814), .CK(n3724), .QN(n925) );
  DFF_X1 reg_r24_q_reg_2_ ( .D(n2813), .CK(n3724), .QN(n926) );
  DFF_X1 reg_r24_q_reg_1_ ( .D(n2812), .CK(n3724), .QN(n927) );
  DFF_X1 reg_r24_q_reg_0_ ( .D(n2811), .CK(n3724), .QN(n928) );
  DFF_X1 reg_r25_q_reg_31_ ( .D(n2810), .CK(n3724), .QN(n929) );
  DFF_X1 reg_r25_q_reg_30_ ( .D(n2809), .CK(n3724), .QN(n930) );
  DFF_X1 reg_r25_q_reg_29_ ( .D(n2808), .CK(n3724), .QN(n931) );
  DFF_X1 reg_r25_q_reg_28_ ( .D(n2807), .CK(n3724), .QN(n932) );
  DFF_X1 reg_r25_q_reg_27_ ( .D(n2806), .CK(n3724), .QN(n933) );
  DFF_X1 reg_r25_q_reg_26_ ( .D(n2805), .CK(n3724), .QN(n934) );
  DFF_X1 reg_r25_q_reg_25_ ( .D(n2804), .CK(n3724), .QN(n935) );
  DFF_X1 reg_r25_q_reg_24_ ( .D(n2803), .CK(n3724), .QN(n936) );
  DFF_X1 reg_r25_q_reg_23_ ( .D(n2802), .CK(n3724), .QN(n937) );
  DFF_X1 reg_r25_q_reg_22_ ( .D(n2801), .CK(n3724), .QN(n938) );
  DFF_X1 reg_r25_q_reg_21_ ( .D(n2800), .CK(n3724), .QN(n939) );
  DFF_X1 reg_r25_q_reg_20_ ( .D(n2799), .CK(n3724), .QN(n940) );
  DFF_X1 reg_r25_q_reg_19_ ( .D(n2798), .CK(n3724), .QN(n941) );
  DFF_X1 reg_r25_q_reg_18_ ( .D(n2797), .CK(n3724), .QN(n942) );
  DFF_X1 reg_r25_q_reg_17_ ( .D(n2796), .CK(n3724), .QN(n943) );
  DFF_X1 reg_r25_q_reg_16_ ( .D(n2795), .CK(n3724), .QN(n944) );
  DFF_X1 reg_r25_q_reg_15_ ( .D(n2794), .CK(n3724), .QN(n945) );
  DFF_X1 reg_r25_q_reg_14_ ( .D(n2793), .CK(n3724), .QN(n946) );
  DFF_X1 reg_r25_q_reg_13_ ( .D(n2792), .CK(n3724), .QN(n947) );
  DFF_X1 reg_r25_q_reg_12_ ( .D(n2791), .CK(n3724), .QN(n948) );
  DFF_X1 reg_r25_q_reg_11_ ( .D(n2790), .CK(n3724), .QN(n949) );
  DFF_X1 reg_r25_q_reg_10_ ( .D(n2789), .CK(n3724), .QN(n950) );
  DFF_X1 reg_r25_q_reg_9_ ( .D(n2788), .CK(n3724), .QN(n951) );
  DFF_X1 reg_r25_q_reg_8_ ( .D(n2787), .CK(n3724), .QN(n952) );
  DFF_X1 reg_r25_q_reg_7_ ( .D(n2786), .CK(n3724), .QN(n953) );
  DFF_X1 reg_r25_q_reg_6_ ( .D(n2785), .CK(n3724), .QN(n954) );
  DFF_X1 reg_r25_q_reg_5_ ( .D(n2784), .CK(n3724), .QN(n955) );
  DFF_X1 reg_r25_q_reg_4_ ( .D(n2783), .CK(n3724), .QN(n956) );
  DFF_X1 reg_r25_q_reg_3_ ( .D(n2782), .CK(n3724), .QN(n957) );
  DFF_X1 reg_r25_q_reg_2_ ( .D(n2781), .CK(n3724), .QN(n958) );
  DFF_X1 reg_r25_q_reg_1_ ( .D(n2780), .CK(n3724), .QN(n959) );
  DFF_X1 reg_r25_q_reg_0_ ( .D(n2779), .CK(n3724), .QN(n960) );
  DFF_X1 reg_r26_q_reg_31_ ( .D(n1009), .CK(n3724), .Q(x26_s10_w[31]) );
  DFF_X1 reg_r26_q_reg_30_ ( .D(n1025), .CK(n3724), .Q(x26_s10_w[30]) );
  DFF_X1 reg_r26_q_reg_29_ ( .D(n1041), .CK(n3724), .Q(x26_s10_w[29]) );
  DFF_X1 reg_r26_q_reg_28_ ( .D(n1057), .CK(n3724), .Q(x26_s10_w[28]) );
  DFF_X1 reg_r26_q_reg_27_ ( .D(n2358), .CK(n3724), .Q(x26_s10_w[27]) );
  DFF_X1 reg_r26_q_reg_26_ ( .D(n3294), .CK(n3724), .Q(x26_s10_w[26]) );
  DFF_X1 reg_r26_q_reg_25_ ( .D(n3310), .CK(n3724), .Q(x26_s10_w[25]) );
  DFF_X1 reg_r26_q_reg_24_ ( .D(n3326), .CK(n3724), .Q(x26_s10_w[24]) );
  DFF_X1 reg_r26_q_reg_23_ ( .D(n3342), .CK(n3724), .Q(x26_s10_w[23]) );
  DFF_X1 reg_r26_q_reg_22_ ( .D(n3358), .CK(n3724), .Q(x26_s10_w[22]) );
  DFF_X1 reg_r26_q_reg_21_ ( .D(n3374), .CK(n3724), .Q(x26_s10_w[21]) );
  DFF_X1 reg_r26_q_reg_20_ ( .D(n3390), .CK(n3724), .Q(x26_s10_w[20]) );
  DFF_X1 reg_r26_q_reg_19_ ( .D(n3406), .CK(n3724), .Q(x26_s10_w[19]) );
  DFF_X1 reg_r26_q_reg_18_ ( .D(n3422), .CK(n3724), .Q(x26_s10_w[18]) );
  DFF_X1 reg_r26_q_reg_17_ ( .D(n3438), .CK(n3724), .Q(x26_s10_w[17]) );
  DFF_X1 reg_r26_q_reg_16_ ( .D(n3454), .CK(n3724), .Q(x26_s10_w[16]) );
  DFF_X1 reg_r26_q_reg_15_ ( .D(n3470), .CK(n3724), .Q(x26_s10_w[15]) );
  DFF_X1 reg_r26_q_reg_14_ ( .D(n3486), .CK(n3724), .Q(x26_s10_w[14]) );
  DFF_X1 reg_r26_q_reg_13_ ( .D(n3502), .CK(n3724), .Q(x26_s10_w[13]) );
  DFF_X1 reg_r26_q_reg_12_ ( .D(n3518), .CK(n3724), .Q(x26_s10_w[12]) );
  DFF_X1 reg_r26_q_reg_11_ ( .D(n3534), .CK(n3724), .Q(x26_s10_w[11]) );
  DFF_X1 reg_r26_q_reg_10_ ( .D(n3550), .CK(n3724), .Q(x26_s10_w[10]) );
  DFF_X1 reg_r26_q_reg_9_ ( .D(n3566), .CK(n3724), .Q(x26_s10_w[9]) );
  DFF_X1 reg_r26_q_reg_8_ ( .D(n3582), .CK(n3724), .Q(x26_s10_w[8]) );
  DFF_X1 reg_r26_q_reg_7_ ( .D(n3598), .CK(n3724), .Q(x26_s10_w[7]) );
  DFF_X1 reg_r26_q_reg_6_ ( .D(n3614), .CK(n3724), .Q(x26_s10_w[6]) );
  DFF_X1 reg_r26_q_reg_5_ ( .D(n3630), .CK(n3724), .Q(x26_s10_w[5]) );
  DFF_X1 reg_r26_q_reg_4_ ( .D(n3646), .CK(n3724), .Q(x26_s10_w[4]) );
  DFF_X1 reg_r26_q_reg_3_ ( .D(n3662), .CK(n3724), .Q(x26_s10_w[3]) );
  DFF_X1 reg_r26_q_reg_2_ ( .D(n3678), .CK(n3724), .Q(x26_s10_w[2]) );
  DFF_X1 reg_r26_q_reg_1_ ( .D(n3694), .CK(n3724), .Q(x26_s10_w[1]) );
  DFF_X1 reg_r26_q_reg_0_ ( .D(n3710), .CK(n3724), .Q(x26_s10_w[0]) );
  NAND4_X1 U2780 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(rd2[9])
         );
  NAND4_X1 U2781 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(rd2[8])
         );
  NAND4_X1 U2782 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(rd2[7])
         );
  NAND4_X1 U2783 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(rd2[6])
         );
  NAND4_X1 U2784 ( .A1(n1169), .A2(n1170), .A3(n1171), .A4(n1172), .ZN(rd2[5])
         );
  NAND4_X1 U2785 ( .A1(n1186), .A2(n1187), .A3(n1188), .A4(n1189), .ZN(rd2[4])
         );
  NAND4_X1 U2786 ( .A1(n1203), .A2(n1204), .A3(n1205), .A4(n1206), .ZN(rd2[3])
         );
  NAND4_X1 U2787 ( .A1(n1220), .A2(n1221), .A3(n1222), .A4(n1223), .ZN(rd2[31]) );
  NAND4_X1 U2788 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(rd2[30]) );
  NAND4_X1 U2789 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(rd2[2])
         );
  NAND4_X1 U2790 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(rd2[29]) );
  NAND4_X1 U2791 ( .A1(n1288), .A2(n1289), .A3(n1290), .A4(n1291), .ZN(rd2[28]) );
  NAND4_X1 U2792 ( .A1(n1305), .A2(n1306), .A3(n1307), .A4(n1308), .ZN(rd2[27]) );
  NAND4_X1 U2793 ( .A1(n1322), .A2(n1323), .A3(n1324), .A4(n1325), .ZN(rd2[26]) );
  NAND4_X1 U2794 ( .A1(n1339), .A2(n1340), .A3(n1341), .A4(n1342), .ZN(rd2[25]) );
  NAND4_X1 U2795 ( .A1(n1356), .A2(n1357), .A3(n1358), .A4(n1359), .ZN(rd2[24]) );
  NAND4_X1 U2796 ( .A1(n1373), .A2(n1374), .A3(n1375), .A4(n1376), .ZN(rd2[23]) );
  NAND4_X1 U2797 ( .A1(n1390), .A2(n1391), .A3(n1392), .A4(n1393), .ZN(rd2[22]) );
  NAND4_X1 U2798 ( .A1(n1407), .A2(n1408), .A3(n1409), .A4(n1410), .ZN(rd2[21]) );
  NAND4_X1 U2799 ( .A1(n1424), .A2(n1425), .A3(n1426), .A4(n1427), .ZN(rd2[20]) );
  NAND4_X1 U2800 ( .A1(n1441), .A2(n1442), .A3(n1443), .A4(n1444), .ZN(rd2[1])
         );
  NAND4_X1 U2801 ( .A1(n1458), .A2(n1459), .A3(n1460), .A4(n1461), .ZN(rd2[19]) );
  NAND4_X1 U2802 ( .A1(n1475), .A2(n1476), .A3(n1477), .A4(n1478), .ZN(rd2[18]) );
  NAND4_X1 U2803 ( .A1(n1492), .A2(n1493), .A3(n1494), .A4(n1495), .ZN(rd2[17]) );
  NAND4_X1 U2804 ( .A1(n1509), .A2(n1510), .A3(n1511), .A4(n1512), .ZN(rd2[16]) );
  NAND4_X1 U2805 ( .A1(n1526), .A2(n1527), .A3(n1528), .A4(n1529), .ZN(rd2[15]) );
  NAND4_X1 U2806 ( .A1(n1543), .A2(n1544), .A3(n1545), .A4(n1546), .ZN(rd2[14]) );
  NAND4_X1 U2807 ( .A1(n1560), .A2(n1561), .A3(n1562), .A4(n1563), .ZN(rd2[13]) );
  NAND4_X1 U2808 ( .A1(n1577), .A2(n1578), .A3(n1579), .A4(n1580), .ZN(rd2[12]) );
  NAND4_X1 U2809 ( .A1(n1594), .A2(n1595), .A3(n1596), .A4(n1597), .ZN(rd2[11]) );
  NAND4_X1 U2810 ( .A1(n1611), .A2(n1612), .A3(n1613), .A4(n1614), .ZN(rd2[10]) );
  NAND4_X1 U2811 ( .A1(n1628), .A2(n1629), .A3(n1630), .A4(n1631), .ZN(rd2[0])
         );
  NAND4_X1 U2812 ( .A1(n1660), .A2(n1661), .A3(n1662), .A4(n1663), .ZN(rd1[9])
         );
  NAND4_X1 U2813 ( .A1(n1708), .A2(n1709), .A3(n1710), .A4(n1711), .ZN(rd1[8])
         );
  NAND4_X1 U2814 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .ZN(rd1[7])
         );
  NAND4_X1 U2815 ( .A1(n1742), .A2(n1743), .A3(n1744), .A4(n1745), .ZN(rd1[6])
         );
  NAND4_X1 U2816 ( .A1(n1759), .A2(n1760), .A3(n1761), .A4(n1762), .ZN(rd1[5])
         );
  NAND4_X1 U2817 ( .A1(n1776), .A2(n1777), .A3(n1778), .A4(n1779), .ZN(rd1[4])
         );
  NAND4_X1 U2818 ( .A1(n1793), .A2(n1794), .A3(n1795), .A4(n1796), .ZN(rd1[3])
         );
  NAND4_X1 U2819 ( .A1(n1810), .A2(n1811), .A3(n1812), .A4(n1813), .ZN(rd1[31]) );
  NAND4_X1 U2820 ( .A1(n1827), .A2(n1828), .A3(n1829), .A4(n1830), .ZN(rd1[30]) );
  NAND4_X1 U2821 ( .A1(n1844), .A2(n1845), .A3(n1846), .A4(n1847), .ZN(rd1[2])
         );
  NAND4_X1 U2822 ( .A1(n1861), .A2(n1862), .A3(n1863), .A4(n1864), .ZN(rd1[29]) );
  NAND4_X1 U2823 ( .A1(n1878), .A2(n1879), .A3(n1880), .A4(n1881), .ZN(rd1[28]) );
  NAND4_X1 U2824 ( .A1(n1895), .A2(n1896), .A3(n1897), .A4(n1898), .ZN(rd1[27]) );
  NAND4_X1 U2825 ( .A1(n1912), .A2(n1913), .A3(n1914), .A4(n1915), .ZN(rd1[26]) );
  NAND4_X1 U2826 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(rd1[25]) );
  NAND4_X1 U2827 ( .A1(n1946), .A2(n1947), .A3(n1948), .A4(n1949), .ZN(rd1[24]) );
  NAND4_X1 U2828 ( .A1(n1963), .A2(n1964), .A3(n1965), .A4(n1966), .ZN(rd1[23]) );
  NAND4_X1 U2829 ( .A1(n1980), .A2(n1981), .A3(n1982), .A4(n1983), .ZN(rd1[22]) );
  NAND4_X1 U2830 ( .A1(n1997), .A2(n1998), .A3(n1999), .A4(n2000), .ZN(rd1[21]) );
  NAND4_X1 U2831 ( .A1(n2014), .A2(n2015), .A3(n2016), .A4(n2017), .ZN(rd1[20]) );
  NAND4_X1 U2832 ( .A1(n2031), .A2(n2032), .A3(n2033), .A4(n2034), .ZN(rd1[1])
         );
  NAND4_X1 U2833 ( .A1(n2048), .A2(n2049), .A3(n2050), .A4(n2051), .ZN(rd1[19]) );
  NAND4_X1 U2834 ( .A1(n2065), .A2(n2066), .A3(n2067), .A4(n2068), .ZN(rd1[18]) );
  NAND4_X1 U2835 ( .A1(n2082), .A2(n2083), .A3(n2084), .A4(n2085), .ZN(rd1[17]) );
  NAND4_X1 U2836 ( .A1(n2099), .A2(n2100), .A3(n2101), .A4(n2102), .ZN(rd1[16]) );
  NAND4_X1 U2837 ( .A1(n2116), .A2(n2117), .A3(n2118), .A4(n2119), .ZN(rd1[15]) );
  NAND4_X1 U2838 ( .A1(n2133), .A2(n2134), .A3(n2135), .A4(n2136), .ZN(rd1[14]) );
  NAND4_X1 U2839 ( .A1(n2150), .A2(n2151), .A3(n2152), .A4(n2153), .ZN(rd1[13]) );
  NAND4_X1 U2840 ( .A1(n2167), .A2(n2168), .A3(n2169), .A4(n2170), .ZN(rd1[12]) );
  NAND4_X1 U2841 ( .A1(n2184), .A2(n2185), .A3(n2186), .A4(n2187), .ZN(rd1[11]) );
  NAND4_X1 U2842 ( .A1(n2201), .A2(n2202), .A3(n2203), .A4(n2204), .ZN(rd1[10]) );
  NAND4_X1 U2843 ( .A1(n2218), .A2(n2219), .A3(n2220), .A4(n2221), .ZN(rd1[0])
         );
  NOR2_X1 U2 ( .A1(n3713), .A2(wa[0]), .ZN(n2283) );
  NOR2_X1 U3 ( .A1(n3714), .A2(n3713), .ZN(n2322) );
  NOR2_X1 U4 ( .A1(n3714), .A2(wa[1]), .ZN(n2286) );
  NOR2_X1 U5 ( .A1(wa[0]), .A2(wa[1]), .ZN(n2288) );
  INV_X1 U6 ( .A(n2290), .ZN(n581) );
  INV_X1 U7 ( .A(n2290), .ZN(n580) );
  INV_X1 U8 ( .A(n2432), .ZN(n381) );
  INV_X1 U9 ( .A(n2432), .ZN(n380) );
  INV_X1 U10 ( .A(n2573), .ZN(n181) );
  INV_X1 U11 ( .A(n2573), .ZN(n180) );
  INV_X1 U12 ( .A(n2678), .ZN(n118) );
  INV_X1 U13 ( .A(n2678), .ZN(n117) );
  INV_X1 U14 ( .A(n2745), .ZN(n100) );
  INV_X1 U15 ( .A(n2745), .ZN(n99) );
  INV_X1 U17 ( .A(n65), .ZN(n416) );
  INV_X1 U19 ( .A(n66), .ZN(n344) );
  INV_X1 U21 ( .A(n67), .ZN(n144) );
  INV_X1 U22 ( .A(n2325), .ZN(n444) );
  INV_X1 U23 ( .A(n2325), .ZN(n443) );
  INV_X1 U24 ( .A(n2365), .ZN(n399) );
  INV_X1 U25 ( .A(n2365), .ZN(n398) );
  INV_X1 U26 ( .A(n2398), .ZN(n390) );
  INV_X1 U27 ( .A(n2398), .ZN(n389) );
  INV_X1 U28 ( .A(n2466), .ZN(n372) );
  INV_X1 U29 ( .A(n2466), .ZN(n371) );
  INV_X1 U30 ( .A(n2506), .ZN(n327) );
  INV_X1 U31 ( .A(n2506), .ZN(n326) );
  INV_X1 U32 ( .A(n2539), .ZN(n190) );
  INV_X1 U33 ( .A(n2539), .ZN(n189) );
  INV_X1 U34 ( .A(n2607), .ZN(n172) );
  INV_X1 U35 ( .A(n2607), .ZN(n171) );
  INV_X1 U36 ( .A(n2645), .ZN(n127) );
  INV_X1 U37 ( .A(n2645), .ZN(n126) );
  INV_X1 U38 ( .A(n2712), .ZN(n109) );
  INV_X1 U39 ( .A(n2712), .ZN(n108) );
  INV_X1 U41 ( .A(n70), .ZN(n598) );
  INV_X1 U43 ( .A(n69), .ZN(n589) );
  INV_X1 U45 ( .A(n71), .ZN(n434) );
  INV_X1 U47 ( .A(n78), .ZN(n425) );
  INV_X1 U49 ( .A(n72), .ZN(n407) );
  INV_X1 U51 ( .A(n73), .ZN(n362) );
  INV_X1 U53 ( .A(n79), .ZN(n353) );
  INV_X1 U55 ( .A(n74), .ZN(n335) );
  INV_X1 U57 ( .A(n75), .ZN(n162) );
  INV_X1 U59 ( .A(n68), .ZN(n153) );
  INV_X1 U61 ( .A(n76), .ZN(n135) );
  INV_X1 U63 ( .A(n77), .ZN(n90) );
  INV_X1 U65 ( .A(n80), .ZN(n81) );
  INV_X1 U66 ( .A(n2251), .ZN(n608) );
  INV_X1 U67 ( .A(n2251), .ZN(n607) );
  AND2_X1 U486 ( .A1(n2360), .A2(n2571), .ZN(n2284) );
  AND2_X1 U492 ( .A1(n2359), .A2(n2360), .ZN(n2323) );
  AND2_X1 U493 ( .A1(n2500), .A2(n2571), .ZN(n2503) );
  AND2_X1 U494 ( .A1(n2500), .A2(n2501), .ZN(n2464) );
  AND2_X1 U495 ( .A1(n2500), .A2(n2359), .ZN(n2605) );
  AND2_X1 U496 ( .A1(n2430), .A2(n2360), .ZN(n2362) );
  AND2_X1 U497 ( .A1(n2501), .A2(n2360), .ZN(n2710) );
  NOR2_X1 U498 ( .A1(n3712), .A2(n3711), .ZN(n2501) );
  AND2_X1 U499 ( .A1(n2500), .A2(n2430), .ZN(n2642) );
  NOR3_X1 U511 ( .A1(n3717), .A2(n3718), .A3(n3716), .ZN(n1648) );
  NOR3_X1 U512 ( .A1(n3721), .A2(n3722), .A3(n3720), .ZN(n2238) );
  AND2_X1 U575 ( .A1(n1656), .A2(n3716), .ZN(n1643) );
  AND2_X1 U576 ( .A1(n1654), .A2(n3717), .ZN(n1640) );
  AND2_X1 U577 ( .A1(n2246), .A2(n3720), .ZN(n2233) );
  AND2_X1 U578 ( .A1(n2244), .A2(n3721), .ZN(n2230) );
  AND2_X1 U579 ( .A1(n1659), .A2(n3718), .ZN(n1646) );
  AND2_X1 U580 ( .A1(n2249), .A2(n3722), .ZN(n2236) );
  INV_X1 U581 ( .A(wdata[0]), .ZN(n3695) );
  INV_X1 U582 ( .A(wdata[1]), .ZN(n3679) );
  INV_X1 U583 ( .A(wdata[2]), .ZN(n3663) );
  INV_X1 U584 ( .A(wdata[3]), .ZN(n3647) );
  INV_X1 U585 ( .A(wdata[4]), .ZN(n3631) );
  INV_X1 U586 ( .A(wdata[5]), .ZN(n3615) );
  INV_X1 U587 ( .A(wdata[6]), .ZN(n3599) );
  INV_X1 U588 ( .A(wdata[7]), .ZN(n3583) );
  INV_X1 U589 ( .A(wdata[8]), .ZN(n3567) );
  INV_X1 U590 ( .A(wdata[9]), .ZN(n3551) );
  INV_X1 U591 ( .A(wdata[10]), .ZN(n3535) );
  INV_X1 U592 ( .A(wdata[11]), .ZN(n3519) );
  INV_X1 U593 ( .A(wdata[12]), .ZN(n3503) );
  INV_X1 U594 ( .A(wdata[13]), .ZN(n3487) );
  INV_X1 U595 ( .A(wdata[14]), .ZN(n3471) );
  INV_X1 U596 ( .A(wdata[15]), .ZN(n3455) );
  INV_X1 U597 ( .A(wdata[16]), .ZN(n3439) );
  INV_X1 U598 ( .A(wdata[17]), .ZN(n3423) );
  INV_X1 U599 ( .A(wdata[18]), .ZN(n3407) );
  INV_X1 U600 ( .A(wdata[19]), .ZN(n3391) );
  INV_X1 U601 ( .A(wdata[20]), .ZN(n3375) );
  INV_X1 U602 ( .A(wdata[21]), .ZN(n3359) );
  INV_X1 U603 ( .A(wdata[22]), .ZN(n3343) );
  INV_X1 U604 ( .A(wdata[23]), .ZN(n3327) );
  INV_X1 U605 ( .A(wdata[24]), .ZN(n3311) );
  INV_X1 U606 ( .A(wdata[25]), .ZN(n3295) );
  INV_X1 U607 ( .A(wdata[26]), .ZN(n2361) );
  INV_X1 U608 ( .A(wdata[27]), .ZN(n1058) );
  INV_X1 U609 ( .A(wdata[28]), .ZN(n1042) );
  INV_X1 U610 ( .A(wdata[29]), .ZN(n1026) );
  INV_X1 U611 ( .A(wdata[30]), .ZN(n1010) );
  INV_X1 U612 ( .A(wdata[31]), .ZN(n994) );
  OAI221_X1 U613 ( .B1(n1078), .B2(n768), .C1(n1079), .C2(n736), .A(n1636), 
        .ZN(n1635) );
  AOI22_X1 U614 ( .A1(x17_a7_w[0]), .A2(n1081), .B1(x16_a6_w[0]), .B2(n1082), 
        .ZN(n1636) );
  OAI221_X1 U615 ( .B1(n1078), .B2(n767), .C1(n1079), .C2(n735), .A(n1449), 
        .ZN(n1448) );
  AOI22_X1 U616 ( .A1(x17_a7_w[1]), .A2(n1081), .B1(x16_a6_w[1]), .B2(n1082), 
        .ZN(n1449) );
  OAI221_X1 U617 ( .B1(n1078), .B2(n766), .C1(n1079), .C2(n734), .A(n1262), 
        .ZN(n1261) );
  AOI22_X1 U618 ( .A1(x17_a7_w[2]), .A2(n1081), .B1(x16_a6_w[2]), .B2(n1082), 
        .ZN(n1262) );
  OAI221_X1 U619 ( .B1(n1078), .B2(n758), .C1(n1079), .C2(n726), .A(n1619), 
        .ZN(n1618) );
  AOI22_X1 U620 ( .A1(x17_a7_w[10]), .A2(n1081), .B1(x16_a6_w[10]), .B2(n1082), 
        .ZN(n1619) );
  OAI221_X1 U621 ( .B1(n1078), .B2(n757), .C1(n1079), .C2(n725), .A(n1602), 
        .ZN(n1601) );
  AOI22_X1 U622 ( .A1(x17_a7_w[11]), .A2(n1081), .B1(x16_a6_w[11]), .B2(n1082), 
        .ZN(n1602) );
  OAI221_X1 U623 ( .B1(n1078), .B2(n756), .C1(n1079), .C2(n724), .A(n1585), 
        .ZN(n1584) );
  AOI22_X1 U624 ( .A1(x17_a7_w[12]), .A2(n1081), .B1(x16_a6_w[12]), .B2(n1082), 
        .ZN(n1585) );
  OAI221_X1 U625 ( .B1(n1078), .B2(n755), .C1(n1079), .C2(n723), .A(n1568), 
        .ZN(n1567) );
  AOI22_X1 U626 ( .A1(x17_a7_w[13]), .A2(n1081), .B1(x16_a6_w[13]), .B2(n1082), 
        .ZN(n1568) );
  OAI221_X1 U627 ( .B1(n1078), .B2(n754), .C1(n1079), .C2(n722), .A(n1551), 
        .ZN(n1550) );
  AOI22_X1 U628 ( .A1(x17_a7_w[14]), .A2(n1081), .B1(x16_a6_w[14]), .B2(n1082), 
        .ZN(n1551) );
  OAI221_X1 U629 ( .B1(n1078), .B2(n753), .C1(n1079), .C2(n721), .A(n1534), 
        .ZN(n1533) );
  AOI22_X1 U630 ( .A1(x17_a7_w[15]), .A2(n1081), .B1(x16_a6_w[15]), .B2(n1082), 
        .ZN(n1534) );
  OAI221_X1 U631 ( .B1(n1078), .B2(n752), .C1(n1079), .C2(n720), .A(n1517), 
        .ZN(n1516) );
  AOI22_X1 U632 ( .A1(x17_a7_w[16]), .A2(n1081), .B1(x16_a6_w[16]), .B2(n1082), 
        .ZN(n1517) );
  OAI221_X1 U633 ( .B1(n1078), .B2(n751), .C1(n1079), .C2(n719), .A(n1500), 
        .ZN(n1499) );
  AOI22_X1 U634 ( .A1(x17_a7_w[17]), .A2(n1081), .B1(x16_a6_w[17]), .B2(n1082), 
        .ZN(n1500) );
  OAI221_X1 U635 ( .B1(n1078), .B2(n750), .C1(n1079), .C2(n718), .A(n1483), 
        .ZN(n1482) );
  AOI22_X1 U636 ( .A1(x17_a7_w[18]), .A2(n1081), .B1(x16_a6_w[18]), .B2(n1082), 
        .ZN(n1483) );
  OAI221_X1 U637 ( .B1(n1078), .B2(n749), .C1(n1079), .C2(n717), .A(n1466), 
        .ZN(n1465) );
  AOI22_X1 U638 ( .A1(x17_a7_w[19]), .A2(n1081), .B1(x16_a6_w[19]), .B2(n1082), 
        .ZN(n1466) );
  OAI221_X1 U639 ( .B1(n1078), .B2(n748), .C1(n1079), .C2(n716), .A(n1432), 
        .ZN(n1431) );
  AOI22_X1 U640 ( .A1(x17_a7_w[20]), .A2(n1081), .B1(x16_a6_w[20]), .B2(n1082), 
        .ZN(n1432) );
  OAI221_X1 U641 ( .B1(n1078), .B2(n747), .C1(n1079), .C2(n715), .A(n1415), 
        .ZN(n1414) );
  AOI22_X1 U642 ( .A1(x17_a7_w[21]), .A2(n1081), .B1(x16_a6_w[21]), .B2(n1082), 
        .ZN(n1415) );
  OAI221_X1 U643 ( .B1(n1078), .B2(n746), .C1(n1079), .C2(n714), .A(n1398), 
        .ZN(n1397) );
  AOI22_X1 U644 ( .A1(x17_a7_w[22]), .A2(n1081), .B1(x16_a6_w[22]), .B2(n1082), 
        .ZN(n1398) );
  OAI221_X1 U645 ( .B1(n1078), .B2(n745), .C1(n1079), .C2(n713), .A(n1381), 
        .ZN(n1380) );
  AOI22_X1 U646 ( .A1(x17_a7_w[23]), .A2(n1081), .B1(x16_a6_w[23]), .B2(n1082), 
        .ZN(n1381) );
  OAI221_X1 U647 ( .B1(n1078), .B2(n744), .C1(n1079), .C2(n712), .A(n1364), 
        .ZN(n1363) );
  AOI22_X1 U648 ( .A1(x17_a7_w[24]), .A2(n1081), .B1(x16_a6_w[24]), .B2(n1082), 
        .ZN(n1364) );
  OAI221_X1 U649 ( .B1(n1078), .B2(n743), .C1(n1079), .C2(n711), .A(n1347), 
        .ZN(n1346) );
  AOI22_X1 U650 ( .A1(x17_a7_w[25]), .A2(n1081), .B1(x16_a6_w[25]), .B2(n1082), 
        .ZN(n1347) );
  OAI221_X1 U651 ( .B1(n1078), .B2(n742), .C1(n1079), .C2(n710), .A(n1330), 
        .ZN(n1329) );
  AOI22_X1 U652 ( .A1(x17_a7_w[26]), .A2(n1081), .B1(x16_a6_w[26]), .B2(n1082), 
        .ZN(n1330) );
  OAI221_X1 U653 ( .B1(n1078), .B2(n741), .C1(n1079), .C2(n709), .A(n1313), 
        .ZN(n1312) );
  AOI22_X1 U654 ( .A1(x17_a7_w[27]), .A2(n1081), .B1(x16_a6_w[27]), .B2(n1082), 
        .ZN(n1313) );
  OAI221_X1 U655 ( .B1(n1078), .B2(n740), .C1(n1079), .C2(n708), .A(n1296), 
        .ZN(n1295) );
  AOI22_X1 U656 ( .A1(x17_a7_w[28]), .A2(n1081), .B1(x16_a6_w[28]), .B2(n1082), 
        .ZN(n1296) );
  OAI221_X1 U657 ( .B1(n1078), .B2(n739), .C1(n1079), .C2(n707), .A(n1279), 
        .ZN(n1278) );
  AOI22_X1 U658 ( .A1(x17_a7_w[29]), .A2(n1081), .B1(x16_a6_w[29]), .B2(n1082), 
        .ZN(n1279) );
  OAI221_X1 U659 ( .B1(n1078), .B2(n738), .C1(n1079), .C2(n706), .A(n1245), 
        .ZN(n1244) );
  AOI22_X1 U660 ( .A1(x17_a7_w[30]), .A2(n1081), .B1(x16_a6_w[30]), .B2(n1082), 
        .ZN(n1245) );
  INV_X1 U661 ( .A(n2406), .ZN(n3578) );
  AOI22_X1 U662 ( .A1(wdata[8]), .A2(n390), .B1(n2398), .B2(x16_a6_w[8]), .ZN(
        n2406) );
  INV_X1 U663 ( .A(n2407), .ZN(n3562) );
  AOI22_X1 U664 ( .A1(wdata[9]), .A2(n390), .B1(n2398), .B2(x16_a6_w[9]), .ZN(
        n2407) );
  INV_X1 U665 ( .A(n2408), .ZN(n3546) );
  AOI22_X1 U666 ( .A1(wdata[10]), .A2(n390), .B1(n2398), .B2(x16_a6_w[10]), 
        .ZN(n2408) );
  INV_X1 U667 ( .A(n2409), .ZN(n3530) );
  AOI22_X1 U668 ( .A1(wdata[11]), .A2(n390), .B1(n2398), .B2(x16_a6_w[11]), 
        .ZN(n2409) );
  INV_X1 U669 ( .A(n2410), .ZN(n3514) );
  AOI22_X1 U670 ( .A1(wdata[12]), .A2(n390), .B1(n2398), .B2(x16_a6_w[12]), 
        .ZN(n2410) );
  INV_X1 U671 ( .A(n2411), .ZN(n3498) );
  AOI22_X1 U672 ( .A1(wdata[13]), .A2(n390), .B1(n2398), .B2(x16_a6_w[13]), 
        .ZN(n2411) );
  INV_X1 U673 ( .A(n2412), .ZN(n3482) );
  AOI22_X1 U674 ( .A1(wdata[14]), .A2(n390), .B1(n2398), .B2(x16_a6_w[14]), 
        .ZN(n2412) );
  INV_X1 U675 ( .A(n2413), .ZN(n3466) );
  AOI22_X1 U676 ( .A1(wdata[15]), .A2(n390), .B1(n2398), .B2(x16_a6_w[15]), 
        .ZN(n2413) );
  INV_X1 U677 ( .A(n2414), .ZN(n3450) );
  AOI22_X1 U678 ( .A1(wdata[16]), .A2(n390), .B1(n2398), .B2(x16_a6_w[16]), 
        .ZN(n2414) );
  INV_X1 U679 ( .A(n2415), .ZN(n3434) );
  AOI22_X1 U680 ( .A1(wdata[17]), .A2(n390), .B1(n2398), .B2(x16_a6_w[17]), 
        .ZN(n2415) );
  INV_X1 U681 ( .A(n2416), .ZN(n3418) );
  AOI22_X1 U682 ( .A1(wdata[18]), .A2(n390), .B1(n2398), .B2(x16_a6_w[18]), 
        .ZN(n2416) );
  INV_X1 U683 ( .A(n2417), .ZN(n3402) );
  AOI22_X1 U684 ( .A1(wdata[19]), .A2(n390), .B1(n2398), .B2(x16_a6_w[19]), 
        .ZN(n2417) );
  INV_X1 U685 ( .A(n2418), .ZN(n3386) );
  AOI22_X1 U686 ( .A1(wdata[20]), .A2(n389), .B1(n2398), .B2(x16_a6_w[20]), 
        .ZN(n2418) );
  INV_X1 U687 ( .A(n2419), .ZN(n3370) );
  AOI22_X1 U688 ( .A1(wdata[21]), .A2(n389), .B1(n2398), .B2(x16_a6_w[21]), 
        .ZN(n2419) );
  INV_X1 U689 ( .A(n2420), .ZN(n3354) );
  AOI22_X1 U690 ( .A1(wdata[22]), .A2(n389), .B1(n2398), .B2(x16_a6_w[22]), 
        .ZN(n2420) );
  INV_X1 U691 ( .A(n2421), .ZN(n3338) );
  AOI22_X1 U692 ( .A1(wdata[23]), .A2(n389), .B1(n2398), .B2(x16_a6_w[23]), 
        .ZN(n2421) );
  INV_X1 U693 ( .A(n2422), .ZN(n3322) );
  AOI22_X1 U694 ( .A1(wdata[24]), .A2(n389), .B1(n2398), .B2(x16_a6_w[24]), 
        .ZN(n2422) );
  INV_X1 U695 ( .A(n2423), .ZN(n3306) );
  AOI22_X1 U696 ( .A1(wdata[25]), .A2(n389), .B1(n2398), .B2(x16_a6_w[25]), 
        .ZN(n2423) );
  INV_X1 U697 ( .A(n2424), .ZN(n2778) );
  AOI22_X1 U698 ( .A1(wdata[26]), .A2(n389), .B1(n2398), .B2(x16_a6_w[26]), 
        .ZN(n2424) );
  INV_X1 U699 ( .A(n2425), .ZN(n1069) );
  AOI22_X1 U700 ( .A1(wdata[27]), .A2(n389), .B1(n2398), .B2(x16_a6_w[27]), 
        .ZN(n2425) );
  INV_X1 U701 ( .A(n2426), .ZN(n1053) );
  AOI22_X1 U702 ( .A1(wdata[28]), .A2(n389), .B1(n2398), .B2(x16_a6_w[28]), 
        .ZN(n2426) );
  INV_X1 U703 ( .A(n2427), .ZN(n1037) );
  AOI22_X1 U704 ( .A1(wdata[29]), .A2(n389), .B1(n2398), .B2(x16_a6_w[29]), 
        .ZN(n2427) );
  INV_X1 U705 ( .A(n2428), .ZN(n1021) );
  AOI22_X1 U706 ( .A1(wdata[30]), .A2(n389), .B1(n2398), .B2(x16_a6_w[30]), 
        .ZN(n2428) );
  INV_X1 U707 ( .A(n2429), .ZN(n1005) );
  AOI22_X1 U708 ( .A1(wdata[31]), .A2(n389), .B1(n2398), .B2(x16_a6_w[31]), 
        .ZN(n2429) );
  OAI221_X1 U709 ( .B1(n1103), .B2(n320), .C1(n1104), .C2(n288), .A(n1655), 
        .ZN(n1650) );
  AOI22_X1 U710 ( .A1(x7_t2_w[0]), .A2(n1106), .B1(x6_t1_w[0]), .B2(n1107), 
        .ZN(n1655) );
  OAI221_X1 U711 ( .B1(n1103), .B2(n319), .C1(n1104), .C2(n287), .A(n1455), 
        .ZN(n1453) );
  AOI22_X1 U712 ( .A1(x7_t2_w[1]), .A2(n1106), .B1(x6_t1_w[1]), .B2(n1107), 
        .ZN(n1455) );
  OAI221_X1 U713 ( .B1(n1103), .B2(n318), .C1(n1104), .C2(n286), .A(n1268), 
        .ZN(n1266) );
  AOI22_X1 U714 ( .A1(x7_t2_w[2]), .A2(n1106), .B1(x6_t1_w[2]), .B2(n1107), 
        .ZN(n1268) );
  OAI221_X1 U715 ( .B1(n1103), .B2(n310), .C1(n1104), .C2(n278), .A(n1625), 
        .ZN(n1623) );
  AOI22_X1 U716 ( .A1(x7_t2_w[10]), .A2(n1106), .B1(x6_t1_w[10]), .B2(n1107), 
        .ZN(n1625) );
  OAI221_X1 U717 ( .B1(n1103), .B2(n309), .C1(n1104), .C2(n277), .A(n1608), 
        .ZN(n1606) );
  AOI22_X1 U718 ( .A1(x7_t2_w[11]), .A2(n1106), .B1(x6_t1_w[11]), .B2(n1107), 
        .ZN(n1608) );
  OAI221_X1 U719 ( .B1(n1103), .B2(n308), .C1(n1104), .C2(n276), .A(n1591), 
        .ZN(n1589) );
  AOI22_X1 U720 ( .A1(x7_t2_w[12]), .A2(n1106), .B1(x6_t1_w[12]), .B2(n1107), 
        .ZN(n1591) );
  OAI221_X1 U721 ( .B1(n1103), .B2(n307), .C1(n1104), .C2(n275), .A(n1574), 
        .ZN(n1572) );
  AOI22_X1 U722 ( .A1(x7_t2_w[13]), .A2(n1106), .B1(x6_t1_w[13]), .B2(n1107), 
        .ZN(n1574) );
  OAI221_X1 U723 ( .B1(n1103), .B2(n306), .C1(n1104), .C2(n274), .A(n1557), 
        .ZN(n1555) );
  AOI22_X1 U724 ( .A1(x7_t2_w[14]), .A2(n1106), .B1(x6_t1_w[14]), .B2(n1107), 
        .ZN(n1557) );
  OAI221_X1 U725 ( .B1(n1103), .B2(n305), .C1(n1104), .C2(n273), .A(n1540), 
        .ZN(n1538) );
  AOI22_X1 U726 ( .A1(x7_t2_w[15]), .A2(n1106), .B1(x6_t1_w[15]), .B2(n1107), 
        .ZN(n1540) );
  OAI221_X1 U727 ( .B1(n1103), .B2(n304), .C1(n1104), .C2(n272), .A(n1523), 
        .ZN(n1521) );
  AOI22_X1 U728 ( .A1(x7_t2_w[16]), .A2(n1106), .B1(x6_t1_w[16]), .B2(n1107), 
        .ZN(n1523) );
  OAI221_X1 U729 ( .B1(n1103), .B2(n303), .C1(n1104), .C2(n271), .A(n1506), 
        .ZN(n1504) );
  AOI22_X1 U730 ( .A1(x7_t2_w[17]), .A2(n1106), .B1(x6_t1_w[17]), .B2(n1107), 
        .ZN(n1506) );
  OAI221_X1 U731 ( .B1(n1103), .B2(n302), .C1(n1104), .C2(n270), .A(n1489), 
        .ZN(n1487) );
  AOI22_X1 U732 ( .A1(x7_t2_w[18]), .A2(n1106), .B1(x6_t1_w[18]), .B2(n1107), 
        .ZN(n1489) );
  OAI221_X1 U733 ( .B1(n1103), .B2(n301), .C1(n1104), .C2(n269), .A(n1472), 
        .ZN(n1470) );
  AOI22_X1 U734 ( .A1(x7_t2_w[19]), .A2(n1106), .B1(x6_t1_w[19]), .B2(n1107), 
        .ZN(n1472) );
  OAI221_X1 U735 ( .B1(n1103), .B2(n300), .C1(n1104), .C2(n268), .A(n1438), 
        .ZN(n1436) );
  AOI22_X1 U736 ( .A1(x7_t2_w[20]), .A2(n1106), .B1(x6_t1_w[20]), .B2(n1107), 
        .ZN(n1438) );
  OAI221_X1 U737 ( .B1(n1103), .B2(n299), .C1(n1104), .C2(n267), .A(n1421), 
        .ZN(n1419) );
  AOI22_X1 U738 ( .A1(x7_t2_w[21]), .A2(n1106), .B1(x6_t1_w[21]), .B2(n1107), 
        .ZN(n1421) );
  OAI221_X1 U739 ( .B1(n1103), .B2(n298), .C1(n1104), .C2(n266), .A(n1404), 
        .ZN(n1402) );
  AOI22_X1 U740 ( .A1(x7_t2_w[22]), .A2(n1106), .B1(x6_t1_w[22]), .B2(n1107), 
        .ZN(n1404) );
  OAI221_X1 U741 ( .B1(n1103), .B2(n297), .C1(n1104), .C2(n265), .A(n1387), 
        .ZN(n1385) );
  AOI22_X1 U742 ( .A1(x7_t2_w[23]), .A2(n1106), .B1(x6_t1_w[23]), .B2(n1107), 
        .ZN(n1387) );
  OAI221_X1 U743 ( .B1(n1103), .B2(n296), .C1(n1104), .C2(n264), .A(n1370), 
        .ZN(n1368) );
  AOI22_X1 U744 ( .A1(x7_t2_w[24]), .A2(n1106), .B1(x6_t1_w[24]), .B2(n1107), 
        .ZN(n1370) );
  OAI221_X1 U745 ( .B1(n1103), .B2(n295), .C1(n1104), .C2(n263), .A(n1353), 
        .ZN(n1351) );
  AOI22_X1 U746 ( .A1(x7_t2_w[25]), .A2(n1106), .B1(x6_t1_w[25]), .B2(n1107), 
        .ZN(n1353) );
  OAI221_X1 U747 ( .B1(n1103), .B2(n294), .C1(n1104), .C2(n262), .A(n1336), 
        .ZN(n1334) );
  AOI22_X1 U748 ( .A1(x7_t2_w[26]), .A2(n1106), .B1(x6_t1_w[26]), .B2(n1107), 
        .ZN(n1336) );
  OAI221_X1 U749 ( .B1(n1103), .B2(n293), .C1(n1104), .C2(n261), .A(n1319), 
        .ZN(n1317) );
  AOI22_X1 U750 ( .A1(x7_t2_w[27]), .A2(n1106), .B1(x6_t1_w[27]), .B2(n1107), 
        .ZN(n1319) );
  OAI221_X1 U751 ( .B1(n1103), .B2(n292), .C1(n1104), .C2(n260), .A(n1302), 
        .ZN(n1300) );
  AOI22_X1 U752 ( .A1(x7_t2_w[28]), .A2(n1106), .B1(x6_t1_w[28]), .B2(n1107), 
        .ZN(n1302) );
  OAI221_X1 U753 ( .B1(n1103), .B2(n291), .C1(n1104), .C2(n259), .A(n1285), 
        .ZN(n1283) );
  AOI22_X1 U754 ( .A1(x7_t2_w[29]), .A2(n1106), .B1(x6_t1_w[29]), .B2(n1107), 
        .ZN(n1285) );
  OAI221_X1 U755 ( .B1(n1103), .B2(n290), .C1(n1104), .C2(n258), .A(n1251), 
        .ZN(n1249) );
  AOI22_X1 U756 ( .A1(x7_t2_w[30]), .A2(n1106), .B1(x6_t1_w[30]), .B2(n1107), 
        .ZN(n1251) );
  NOR4_X1 U757 ( .A1(n1632), .A2(n1633), .A3(n1634), .A4(n1635), .ZN(n1631) );
  OAI221_X1 U758 ( .B1(n1093), .B2(n64), .C1(n1094), .C2(n32), .A(n1647), .ZN(
        n1632) );
  OAI221_X1 U759 ( .B1(n1088), .B2(n960), .C1(n1089), .C2(n928), .A(n1644), 
        .ZN(n1633) );
  OAI221_X1 U760 ( .B1(n1083), .B2(n832), .C1(n1084), .C2(n800), .A(n1641), 
        .ZN(n1634) );
  NOR4_X1 U761 ( .A1(n1445), .A2(n1446), .A3(n1447), .A4(n1448), .ZN(n1444) );
  OAI221_X1 U762 ( .B1(n1093), .B2(n63), .C1(n1094), .C2(n31), .A(n1452), .ZN(
        n1445) );
  OAI221_X1 U763 ( .B1(n1088), .B2(n959), .C1(n1089), .C2(n927), .A(n1451), 
        .ZN(n1446) );
  OAI221_X1 U764 ( .B1(n1083), .B2(n831), .C1(n1084), .C2(n799), .A(n1450), 
        .ZN(n1447) );
  NOR4_X1 U765 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1257) );
  OAI221_X1 U766 ( .B1(n1093), .B2(n62), .C1(n1094), .C2(n30), .A(n1265), .ZN(
        n1258) );
  OAI221_X1 U767 ( .B1(n1088), .B2(n958), .C1(n1089), .C2(n926), .A(n1264), 
        .ZN(n1259) );
  OAI221_X1 U768 ( .B1(n1083), .B2(n830), .C1(n1084), .C2(n798), .A(n1263), 
        .ZN(n1260) );
  NOR4_X1 U769 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206) );
  OAI221_X1 U770 ( .B1(n1093), .B2(n61), .C1(n1094), .C2(n29), .A(n1214), .ZN(
        n1207) );
  OAI221_X1 U771 ( .B1(n1088), .B2(n957), .C1(n1089), .C2(n925), .A(n1213), 
        .ZN(n1208) );
  OAI221_X1 U772 ( .B1(n1083), .B2(n829), .C1(n1084), .C2(n797), .A(n1212), 
        .ZN(n1209) );
  NOR4_X1 U773 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
  OAI221_X1 U774 ( .B1(n1093), .B2(n60), .C1(n1094), .C2(n28), .A(n1197), .ZN(
        n1190) );
  OAI221_X1 U775 ( .B1(n1088), .B2(n956), .C1(n1089), .C2(n924), .A(n1196), 
        .ZN(n1191) );
  OAI221_X1 U776 ( .B1(n1083), .B2(n828), .C1(n1084), .C2(n796), .A(n1195), 
        .ZN(n1192) );
  NOR4_X1 U777 ( .A1(n1173), .A2(n1174), .A3(n1175), .A4(n1176), .ZN(n1172) );
  OAI221_X1 U778 ( .B1(n1093), .B2(n59), .C1(n1094), .C2(n27), .A(n1180), .ZN(
        n1173) );
  OAI221_X1 U779 ( .B1(n1088), .B2(n955), .C1(n1089), .C2(n923), .A(n1179), 
        .ZN(n1174) );
  OAI221_X1 U780 ( .B1(n1083), .B2(n827), .C1(n1084), .C2(n795), .A(n1178), 
        .ZN(n1175) );
  NOR4_X1 U781 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
  OAI221_X1 U782 ( .B1(n1093), .B2(n58), .C1(n1094), .C2(n26), .A(n1163), .ZN(
        n1156) );
  OAI221_X1 U783 ( .B1(n1088), .B2(n954), .C1(n1089), .C2(n922), .A(n1162), 
        .ZN(n1157) );
  OAI221_X1 U784 ( .B1(n1083), .B2(n826), .C1(n1084), .C2(n794), .A(n1161), 
        .ZN(n1158) );
  NOR4_X1 U785 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1138) );
  OAI221_X1 U786 ( .B1(n1093), .B2(n57), .C1(n1094), .C2(n25), .A(n1146), .ZN(
        n1139) );
  OAI221_X1 U787 ( .B1(n1088), .B2(n953), .C1(n1089), .C2(n921), .A(n1145), 
        .ZN(n1140) );
  OAI221_X1 U788 ( .B1(n1083), .B2(n825), .C1(n1084), .C2(n793), .A(n1144), 
        .ZN(n1141) );
  NOR4_X1 U789 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1121) );
  OAI221_X1 U790 ( .B1(n1093), .B2(n56), .C1(n1094), .C2(n24), .A(n1129), .ZN(
        n1122) );
  OAI221_X1 U791 ( .B1(n1088), .B2(n952), .C1(n1089), .C2(n920), .A(n1128), 
        .ZN(n1123) );
  OAI221_X1 U792 ( .B1(n1083), .B2(n824), .C1(n1084), .C2(n792), .A(n1127), 
        .ZN(n1124) );
  NOR4_X1 U793 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073) );
  OAI221_X1 U794 ( .B1(n1093), .B2(n55), .C1(n1094), .C2(n23), .A(n1095), .ZN(
        n1074) );
  OAI221_X1 U795 ( .B1(n1088), .B2(n951), .C1(n1089), .C2(n919), .A(n1090), 
        .ZN(n1075) );
  OAI221_X1 U796 ( .B1(n1083), .B2(n823), .C1(n1084), .C2(n791), .A(n1085), 
        .ZN(n1076) );
  NOR4_X1 U797 ( .A1(n1615), .A2(n1616), .A3(n1617), .A4(n1618), .ZN(n1614) );
  OAI221_X1 U798 ( .B1(n1093), .B2(n54), .C1(n1094), .C2(n22), .A(n1622), .ZN(
        n1615) );
  OAI221_X1 U799 ( .B1(n1088), .B2(n950), .C1(n1089), .C2(n918), .A(n1621), 
        .ZN(n1616) );
  OAI221_X1 U800 ( .B1(n1083), .B2(n822), .C1(n1084), .C2(n790), .A(n1620), 
        .ZN(n1617) );
  NOR4_X1 U801 ( .A1(n1598), .A2(n1599), .A3(n1600), .A4(n1601), .ZN(n1597) );
  OAI221_X1 U802 ( .B1(n1093), .B2(n53), .C1(n1094), .C2(n21), .A(n1605), .ZN(
        n1598) );
  OAI221_X1 U803 ( .B1(n1088), .B2(n949), .C1(n1089), .C2(n917), .A(n1604), 
        .ZN(n1599) );
  OAI221_X1 U804 ( .B1(n1083), .B2(n821), .C1(n1084), .C2(n789), .A(n1603), 
        .ZN(n1600) );
  NOR4_X1 U805 ( .A1(n1581), .A2(n1582), .A3(n1583), .A4(n1584), .ZN(n1580) );
  OAI221_X1 U806 ( .B1(n1093), .B2(n52), .C1(n1094), .C2(n20), .A(n1588), .ZN(
        n1581) );
  OAI221_X1 U807 ( .B1(n1088), .B2(n948), .C1(n1089), .C2(n916), .A(n1587), 
        .ZN(n1582) );
  OAI221_X1 U808 ( .B1(n1083), .B2(n820), .C1(n1084), .C2(n788), .A(n1586), 
        .ZN(n1583) );
  NOR4_X1 U809 ( .A1(n1564), .A2(n1565), .A3(n1566), .A4(n1567), .ZN(n1563) );
  OAI221_X1 U810 ( .B1(n1093), .B2(n51), .C1(n1094), .C2(n19), .A(n1571), .ZN(
        n1564) );
  OAI221_X1 U811 ( .B1(n1088), .B2(n947), .C1(n1089), .C2(n915), .A(n1570), 
        .ZN(n1565) );
  OAI221_X1 U812 ( .B1(n1083), .B2(n819), .C1(n1084), .C2(n787), .A(n1569), 
        .ZN(n1566) );
  NOR4_X1 U813 ( .A1(n1547), .A2(n1548), .A3(n1549), .A4(n1550), .ZN(n1546) );
  OAI221_X1 U814 ( .B1(n1093), .B2(n50), .C1(n1094), .C2(n18), .A(n1554), .ZN(
        n1547) );
  OAI221_X1 U815 ( .B1(n1088), .B2(n946), .C1(n1089), .C2(n914), .A(n1553), 
        .ZN(n1548) );
  OAI221_X1 U816 ( .B1(n1083), .B2(n818), .C1(n1084), .C2(n786), .A(n1552), 
        .ZN(n1549) );
  NOR4_X1 U817 ( .A1(n1530), .A2(n1531), .A3(n1532), .A4(n1533), .ZN(n1529) );
  OAI221_X1 U818 ( .B1(n1093), .B2(n49), .C1(n1094), .C2(n17), .A(n1537), .ZN(
        n1530) );
  OAI221_X1 U819 ( .B1(n1088), .B2(n945), .C1(n1089), .C2(n913), .A(n1536), 
        .ZN(n1531) );
  OAI221_X1 U820 ( .B1(n1083), .B2(n817), .C1(n1084), .C2(n785), .A(n1535), 
        .ZN(n1532) );
  NOR4_X1 U821 ( .A1(n1513), .A2(n1514), .A3(n1515), .A4(n1516), .ZN(n1512) );
  OAI221_X1 U822 ( .B1(n1093), .B2(n48), .C1(n1094), .C2(n16), .A(n1520), .ZN(
        n1513) );
  OAI221_X1 U823 ( .B1(n1088), .B2(n944), .C1(n1089), .C2(n912), .A(n1519), 
        .ZN(n1514) );
  OAI221_X1 U824 ( .B1(n1083), .B2(n816), .C1(n1084), .C2(n784), .A(n1518), 
        .ZN(n1515) );
  NOR4_X1 U825 ( .A1(n1496), .A2(n1497), .A3(n1498), .A4(n1499), .ZN(n1495) );
  OAI221_X1 U826 ( .B1(n1093), .B2(n47), .C1(n1094), .C2(n15), .A(n1503), .ZN(
        n1496) );
  OAI221_X1 U827 ( .B1(n1088), .B2(n943), .C1(n1089), .C2(n911), .A(n1502), 
        .ZN(n1497) );
  OAI221_X1 U828 ( .B1(n1083), .B2(n815), .C1(n1084), .C2(n783), .A(n1501), 
        .ZN(n1498) );
  NOR4_X1 U829 ( .A1(n1479), .A2(n1480), .A3(n1481), .A4(n1482), .ZN(n1478) );
  OAI221_X1 U830 ( .B1(n1093), .B2(n46), .C1(n1094), .C2(n14), .A(n1486), .ZN(
        n1479) );
  OAI221_X1 U831 ( .B1(n1088), .B2(n942), .C1(n1089), .C2(n910), .A(n1485), 
        .ZN(n1480) );
  OAI221_X1 U832 ( .B1(n1083), .B2(n814), .C1(n1084), .C2(n782), .A(n1484), 
        .ZN(n1481) );
  NOR4_X1 U833 ( .A1(n1462), .A2(n1463), .A3(n1464), .A4(n1465), .ZN(n1461) );
  OAI221_X1 U834 ( .B1(n1093), .B2(n45), .C1(n1094), .C2(n13), .A(n1469), .ZN(
        n1462) );
  OAI221_X1 U835 ( .B1(n1088), .B2(n941), .C1(n1089), .C2(n909), .A(n1468), 
        .ZN(n1463) );
  OAI221_X1 U836 ( .B1(n1083), .B2(n813), .C1(n1084), .C2(n781), .A(n1467), 
        .ZN(n1464) );
  NOR4_X1 U837 ( .A1(n1428), .A2(n1429), .A3(n1430), .A4(n1431), .ZN(n1427) );
  OAI221_X1 U838 ( .B1(n1093), .B2(n44), .C1(n1094), .C2(n12), .A(n1435), .ZN(
        n1428) );
  OAI221_X1 U839 ( .B1(n1088), .B2(n940), .C1(n1089), .C2(n908), .A(n1434), 
        .ZN(n1429) );
  OAI221_X1 U840 ( .B1(n1083), .B2(n812), .C1(n1084), .C2(n780), .A(n1433), 
        .ZN(n1430) );
  NOR4_X1 U841 ( .A1(n1411), .A2(n1412), .A3(n1413), .A4(n1414), .ZN(n1410) );
  OAI221_X1 U842 ( .B1(n1093), .B2(n43), .C1(n1094), .C2(n11), .A(n1418), .ZN(
        n1411) );
  OAI221_X1 U843 ( .B1(n1088), .B2(n939), .C1(n1089), .C2(n907), .A(n1417), 
        .ZN(n1412) );
  OAI221_X1 U844 ( .B1(n1083), .B2(n811), .C1(n1084), .C2(n779), .A(n1416), 
        .ZN(n1413) );
  NOR4_X1 U845 ( .A1(n1394), .A2(n1395), .A3(n1396), .A4(n1397), .ZN(n1393) );
  OAI221_X1 U846 ( .B1(n1093), .B2(n42), .C1(n1094), .C2(n10), .A(n1401), .ZN(
        n1394) );
  OAI221_X1 U847 ( .B1(n1088), .B2(n938), .C1(n1089), .C2(n906), .A(n1400), 
        .ZN(n1395) );
  OAI221_X1 U848 ( .B1(n1083), .B2(n810), .C1(n1084), .C2(n778), .A(n1399), 
        .ZN(n1396) );
  NOR4_X1 U849 ( .A1(n1377), .A2(n1378), .A3(n1379), .A4(n1380), .ZN(n1376) );
  OAI221_X1 U850 ( .B1(n1093), .B2(n41), .C1(n1094), .C2(n9), .A(n1384), .ZN(
        n1377) );
  OAI221_X1 U851 ( .B1(n1088), .B2(n937), .C1(n1089), .C2(n905), .A(n1383), 
        .ZN(n1378) );
  OAI221_X1 U852 ( .B1(n1083), .B2(n809), .C1(n1084), .C2(n777), .A(n1382), 
        .ZN(n1379) );
  NOR4_X1 U853 ( .A1(n1360), .A2(n1361), .A3(n1362), .A4(n1363), .ZN(n1359) );
  OAI221_X1 U854 ( .B1(n1093), .B2(n40), .C1(n1094), .C2(n8), .A(n1367), .ZN(
        n1360) );
  OAI221_X1 U855 ( .B1(n1088), .B2(n936), .C1(n1089), .C2(n904), .A(n1366), 
        .ZN(n1361) );
  OAI221_X1 U856 ( .B1(n1083), .B2(n808), .C1(n1084), .C2(n776), .A(n1365), 
        .ZN(n1362) );
  NOR4_X1 U857 ( .A1(n1343), .A2(n1344), .A3(n1345), .A4(n1346), .ZN(n1342) );
  OAI221_X1 U858 ( .B1(n1093), .B2(n39), .C1(n1094), .C2(n7), .A(n1350), .ZN(
        n1343) );
  OAI221_X1 U859 ( .B1(n1088), .B2(n935), .C1(n1089), .C2(n903), .A(n1349), 
        .ZN(n1344) );
  OAI221_X1 U860 ( .B1(n1083), .B2(n807), .C1(n1084), .C2(n775), .A(n1348), 
        .ZN(n1345) );
  NOR4_X1 U861 ( .A1(n1326), .A2(n1327), .A3(n1328), .A4(n1329), .ZN(n1325) );
  OAI221_X1 U862 ( .B1(n1093), .B2(n38), .C1(n1094), .C2(n6), .A(n1333), .ZN(
        n1326) );
  OAI221_X1 U863 ( .B1(n1088), .B2(n934), .C1(n1089), .C2(n902), .A(n1332), 
        .ZN(n1327) );
  OAI221_X1 U864 ( .B1(n1083), .B2(n806), .C1(n1084), .C2(n774), .A(n1331), 
        .ZN(n1328) );
  NOR4_X1 U865 ( .A1(n1309), .A2(n1310), .A3(n1311), .A4(n1312), .ZN(n1308) );
  OAI221_X1 U866 ( .B1(n1093), .B2(n37), .C1(n1094), .C2(n5), .A(n1316), .ZN(
        n1309) );
  OAI221_X1 U867 ( .B1(n1088), .B2(n933), .C1(n1089), .C2(n901), .A(n1315), 
        .ZN(n1310) );
  OAI221_X1 U868 ( .B1(n1083), .B2(n805), .C1(n1084), .C2(n773), .A(n1314), 
        .ZN(n1311) );
  NOR4_X1 U869 ( .A1(n1292), .A2(n1293), .A3(n1294), .A4(n1295), .ZN(n1291) );
  OAI221_X1 U870 ( .B1(n1093), .B2(n36), .C1(n1094), .C2(n4), .A(n1299), .ZN(
        n1292) );
  OAI221_X1 U871 ( .B1(n1088), .B2(n932), .C1(n1089), .C2(n900), .A(n1298), 
        .ZN(n1293) );
  OAI221_X1 U872 ( .B1(n1083), .B2(n804), .C1(n1084), .C2(n772), .A(n1297), 
        .ZN(n1294) );
  NOR4_X1 U873 ( .A1(n1275), .A2(n1276), .A3(n1277), .A4(n1278), .ZN(n1274) );
  OAI221_X1 U874 ( .B1(n1093), .B2(n35), .C1(n1094), .C2(n3), .A(n1282), .ZN(
        n1275) );
  OAI221_X1 U875 ( .B1(n1088), .B2(n931), .C1(n1089), .C2(n899), .A(n1281), 
        .ZN(n1276) );
  OAI221_X1 U876 ( .B1(n1083), .B2(n803), .C1(n1084), .C2(n771), .A(n1280), 
        .ZN(n1277) );
  NOR4_X1 U877 ( .A1(n1241), .A2(n1242), .A3(n1243), .A4(n1244), .ZN(n1240) );
  OAI221_X1 U878 ( .B1(n1093), .B2(n34), .C1(n1094), .C2(n2), .A(n1248), .ZN(
        n1241) );
  OAI221_X1 U879 ( .B1(n1088), .B2(n930), .C1(n1089), .C2(n898), .A(n1247), 
        .ZN(n1242) );
  OAI221_X1 U880 ( .B1(n1083), .B2(n802), .C1(n1084), .C2(n770), .A(n1246), 
        .ZN(n1243) );
  NOR4_X1 U881 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
  OAI221_X1 U882 ( .B1(n1093), .B2(n33), .C1(n1094), .C2(n1), .A(n1231), .ZN(
        n1224) );
  OAI221_X1 U883 ( .B1(n1088), .B2(n929), .C1(n1089), .C2(n897), .A(n1230), 
        .ZN(n1225) );
  OAI221_X1 U884 ( .B1(n1083), .B2(n801), .C1(n1084), .C2(n769), .A(n1229), 
        .ZN(n1226) );
  NOR4_X1 U885 ( .A1(n2222), .A2(n2223), .A3(n2224), .A4(n2225), .ZN(n2221) );
  OAI221_X1 U886 ( .B1(n64), .B2(n1683), .C1(n32), .C2(n1684), .A(n2237), .ZN(
        n2222) );
  OAI221_X1 U887 ( .B1(n960), .B2(n1678), .C1(n928), .C2(n1679), .A(n2234), 
        .ZN(n2223) );
  OAI221_X1 U888 ( .B1(n832), .B2(n1673), .C1(n800), .C2(n1674), .A(n2231), 
        .ZN(n2224) );
  NOR4_X1 U889 ( .A1(n2035), .A2(n2036), .A3(n2037), .A4(n2038), .ZN(n2034) );
  OAI221_X1 U890 ( .B1(n63), .B2(n1683), .C1(n31), .C2(n1684), .A(n2042), .ZN(
        n2035) );
  OAI221_X1 U891 ( .B1(n959), .B2(n1678), .C1(n927), .C2(n1679), .A(n2041), 
        .ZN(n2036) );
  OAI221_X1 U892 ( .B1(n831), .B2(n1673), .C1(n799), .C2(n1674), .A(n2040), 
        .ZN(n2037) );
  NOR4_X1 U893 ( .A1(n1848), .A2(n1849), .A3(n1850), .A4(n1851), .ZN(n1847) );
  OAI221_X1 U894 ( .B1(n62), .B2(n1683), .C1(n30), .C2(n1684), .A(n1855), .ZN(
        n1848) );
  OAI221_X1 U895 ( .B1(n958), .B2(n1678), .C1(n926), .C2(n1679), .A(n1854), 
        .ZN(n1849) );
  OAI221_X1 U896 ( .B1(n830), .B2(n1673), .C1(n798), .C2(n1674), .A(n1853), 
        .ZN(n1850) );
  NOR4_X1 U897 ( .A1(n1797), .A2(n1798), .A3(n1799), .A4(n1800), .ZN(n1796) );
  OAI221_X1 U898 ( .B1(n61), .B2(n1683), .C1(n29), .C2(n1684), .A(n1804), .ZN(
        n1797) );
  OAI221_X1 U899 ( .B1(n957), .B2(n1678), .C1(n925), .C2(n1679), .A(n1803), 
        .ZN(n1798) );
  OAI221_X1 U900 ( .B1(n829), .B2(n1673), .C1(n797), .C2(n1674), .A(n1802), 
        .ZN(n1799) );
  NOR4_X1 U901 ( .A1(n1780), .A2(n1781), .A3(n1782), .A4(n1783), .ZN(n1779) );
  OAI221_X1 U902 ( .B1(n60), .B2(n1683), .C1(n28), .C2(n1684), .A(n1787), .ZN(
        n1780) );
  OAI221_X1 U903 ( .B1(n956), .B2(n1678), .C1(n924), .C2(n1679), .A(n1786), 
        .ZN(n1781) );
  OAI221_X1 U904 ( .B1(n828), .B2(n1673), .C1(n796), .C2(n1674), .A(n1785), 
        .ZN(n1782) );
  NOR4_X1 U905 ( .A1(n1763), .A2(n1764), .A3(n1765), .A4(n1766), .ZN(n1762) );
  OAI221_X1 U906 ( .B1(n59), .B2(n1683), .C1(n27), .C2(n1684), .A(n1770), .ZN(
        n1763) );
  OAI221_X1 U907 ( .B1(n955), .B2(n1678), .C1(n923), .C2(n1679), .A(n1769), 
        .ZN(n1764) );
  OAI221_X1 U908 ( .B1(n827), .B2(n1673), .C1(n795), .C2(n1674), .A(n1768), 
        .ZN(n1765) );
  NOR4_X1 U909 ( .A1(n1746), .A2(n1747), .A3(n1748), .A4(n1749), .ZN(n1745) );
  OAI221_X1 U910 ( .B1(n58), .B2(n1683), .C1(n26), .C2(n1684), .A(n1753), .ZN(
        n1746) );
  OAI221_X1 U911 ( .B1(n954), .B2(n1678), .C1(n922), .C2(n1679), .A(n1752), 
        .ZN(n1747) );
  OAI221_X1 U912 ( .B1(n826), .B2(n1673), .C1(n794), .C2(n1674), .A(n1751), 
        .ZN(n1748) );
  NOR4_X1 U913 ( .A1(n1729), .A2(n1730), .A3(n1731), .A4(n1732), .ZN(n1728) );
  OAI221_X1 U914 ( .B1(n57), .B2(n1683), .C1(n25), .C2(n1684), .A(n1736), .ZN(
        n1729) );
  OAI221_X1 U915 ( .B1(n953), .B2(n1678), .C1(n921), .C2(n1679), .A(n1735), 
        .ZN(n1730) );
  OAI221_X1 U916 ( .B1(n825), .B2(n1673), .C1(n793), .C2(n1674), .A(n1734), 
        .ZN(n1731) );
  NOR4_X1 U917 ( .A1(n1712), .A2(n1713), .A3(n1714), .A4(n1715), .ZN(n1711) );
  OAI221_X1 U918 ( .B1(n56), .B2(n1683), .C1(n24), .C2(n1684), .A(n1719), .ZN(
        n1712) );
  OAI221_X1 U919 ( .B1(n952), .B2(n1678), .C1(n920), .C2(n1679), .A(n1718), 
        .ZN(n1713) );
  OAI221_X1 U920 ( .B1(n824), .B2(n1673), .C1(n792), .C2(n1674), .A(n1717), 
        .ZN(n1714) );
  NOR4_X1 U921 ( .A1(n1664), .A2(n1665), .A3(n1666), .A4(n1667), .ZN(n1663) );
  OAI221_X1 U922 ( .B1(n55), .B2(n1683), .C1(n23), .C2(n1684), .A(n1685), .ZN(
        n1664) );
  OAI221_X1 U923 ( .B1(n951), .B2(n1678), .C1(n919), .C2(n1679), .A(n1680), 
        .ZN(n1665) );
  OAI221_X1 U924 ( .B1(n823), .B2(n1673), .C1(n791), .C2(n1674), .A(n1675), 
        .ZN(n1666) );
  NOR4_X1 U925 ( .A1(n2205), .A2(n2206), .A3(n2207), .A4(n2208), .ZN(n2204) );
  OAI221_X1 U926 ( .B1(n54), .B2(n1683), .C1(n22), .C2(n1684), .A(n2212), .ZN(
        n2205) );
  OAI221_X1 U927 ( .B1(n950), .B2(n1678), .C1(n918), .C2(n1679), .A(n2211), 
        .ZN(n2206) );
  OAI221_X1 U928 ( .B1(n822), .B2(n1673), .C1(n790), .C2(n1674), .A(n2210), 
        .ZN(n2207) );
  NOR4_X1 U929 ( .A1(n2188), .A2(n2189), .A3(n2190), .A4(n2191), .ZN(n2187) );
  OAI221_X1 U930 ( .B1(n53), .B2(n1683), .C1(n21), .C2(n1684), .A(n2195), .ZN(
        n2188) );
  OAI221_X1 U931 ( .B1(n949), .B2(n1678), .C1(n917), .C2(n1679), .A(n2194), 
        .ZN(n2189) );
  OAI221_X1 U932 ( .B1(n821), .B2(n1673), .C1(n789), .C2(n1674), .A(n2193), 
        .ZN(n2190) );
  NOR4_X1 U933 ( .A1(n2171), .A2(n2172), .A3(n2173), .A4(n2174), .ZN(n2170) );
  OAI221_X1 U934 ( .B1(n52), .B2(n1683), .C1(n20), .C2(n1684), .A(n2178), .ZN(
        n2171) );
  OAI221_X1 U935 ( .B1(n948), .B2(n1678), .C1(n916), .C2(n1679), .A(n2177), 
        .ZN(n2172) );
  OAI221_X1 U936 ( .B1(n820), .B2(n1673), .C1(n788), .C2(n1674), .A(n2176), 
        .ZN(n2173) );
  NOR4_X1 U937 ( .A1(n2154), .A2(n2155), .A3(n2156), .A4(n2157), .ZN(n2153) );
  OAI221_X1 U938 ( .B1(n51), .B2(n1683), .C1(n19), .C2(n1684), .A(n2161), .ZN(
        n2154) );
  OAI221_X1 U939 ( .B1(n947), .B2(n1678), .C1(n915), .C2(n1679), .A(n2160), 
        .ZN(n2155) );
  OAI221_X1 U940 ( .B1(n819), .B2(n1673), .C1(n787), .C2(n1674), .A(n2159), 
        .ZN(n2156) );
  NOR4_X1 U941 ( .A1(n2137), .A2(n2138), .A3(n2139), .A4(n2140), .ZN(n2136) );
  OAI221_X1 U942 ( .B1(n50), .B2(n1683), .C1(n18), .C2(n1684), .A(n2144), .ZN(
        n2137) );
  OAI221_X1 U943 ( .B1(n946), .B2(n1678), .C1(n914), .C2(n1679), .A(n2143), 
        .ZN(n2138) );
  OAI221_X1 U944 ( .B1(n818), .B2(n1673), .C1(n786), .C2(n1674), .A(n2142), 
        .ZN(n2139) );
  NOR4_X1 U945 ( .A1(n2120), .A2(n2121), .A3(n2122), .A4(n2123), .ZN(n2119) );
  OAI221_X1 U946 ( .B1(n49), .B2(n1683), .C1(n17), .C2(n1684), .A(n2127), .ZN(
        n2120) );
  OAI221_X1 U947 ( .B1(n945), .B2(n1678), .C1(n913), .C2(n1679), .A(n2126), 
        .ZN(n2121) );
  OAI221_X1 U948 ( .B1(n817), .B2(n1673), .C1(n785), .C2(n1674), .A(n2125), 
        .ZN(n2122) );
  NOR4_X1 U949 ( .A1(n2103), .A2(n2104), .A3(n2105), .A4(n2106), .ZN(n2102) );
  OAI221_X1 U950 ( .B1(n48), .B2(n1683), .C1(n16), .C2(n1684), .A(n2110), .ZN(
        n2103) );
  OAI221_X1 U951 ( .B1(n944), .B2(n1678), .C1(n912), .C2(n1679), .A(n2109), 
        .ZN(n2104) );
  OAI221_X1 U952 ( .B1(n816), .B2(n1673), .C1(n784), .C2(n1674), .A(n2108), 
        .ZN(n2105) );
  NOR4_X1 U953 ( .A1(n2086), .A2(n2087), .A3(n2088), .A4(n2089), .ZN(n2085) );
  OAI221_X1 U954 ( .B1(n47), .B2(n1683), .C1(n15), .C2(n1684), .A(n2093), .ZN(
        n2086) );
  OAI221_X1 U955 ( .B1(n943), .B2(n1678), .C1(n911), .C2(n1679), .A(n2092), 
        .ZN(n2087) );
  OAI221_X1 U956 ( .B1(n815), .B2(n1673), .C1(n783), .C2(n1674), .A(n2091), 
        .ZN(n2088) );
  NOR4_X1 U957 ( .A1(n2069), .A2(n2070), .A3(n2071), .A4(n2072), .ZN(n2068) );
  OAI221_X1 U958 ( .B1(n46), .B2(n1683), .C1(n14), .C2(n1684), .A(n2076), .ZN(
        n2069) );
  OAI221_X1 U959 ( .B1(n942), .B2(n1678), .C1(n910), .C2(n1679), .A(n2075), 
        .ZN(n2070) );
  OAI221_X1 U960 ( .B1(n814), .B2(n1673), .C1(n782), .C2(n1674), .A(n2074), 
        .ZN(n2071) );
  NOR4_X1 U961 ( .A1(n2052), .A2(n2053), .A3(n2054), .A4(n2055), .ZN(n2051) );
  OAI221_X1 U962 ( .B1(n45), .B2(n1683), .C1(n13), .C2(n1684), .A(n2059), .ZN(
        n2052) );
  OAI221_X1 U963 ( .B1(n941), .B2(n1678), .C1(n909), .C2(n1679), .A(n2058), 
        .ZN(n2053) );
  OAI221_X1 U964 ( .B1(n813), .B2(n1673), .C1(n781), .C2(n1674), .A(n2057), 
        .ZN(n2054) );
  NOR4_X1 U965 ( .A1(n2018), .A2(n2019), .A3(n2020), .A4(n2021), .ZN(n2017) );
  OAI221_X1 U966 ( .B1(n44), .B2(n1683), .C1(n12), .C2(n1684), .A(n2025), .ZN(
        n2018) );
  OAI221_X1 U967 ( .B1(n940), .B2(n1678), .C1(n908), .C2(n1679), .A(n2024), 
        .ZN(n2019) );
  OAI221_X1 U968 ( .B1(n812), .B2(n1673), .C1(n780), .C2(n1674), .A(n2023), 
        .ZN(n2020) );
  NOR4_X1 U969 ( .A1(n2001), .A2(n2002), .A3(n2003), .A4(n2004), .ZN(n2000) );
  OAI221_X1 U970 ( .B1(n43), .B2(n1683), .C1(n11), .C2(n1684), .A(n2008), .ZN(
        n2001) );
  OAI221_X1 U971 ( .B1(n939), .B2(n1678), .C1(n907), .C2(n1679), .A(n2007), 
        .ZN(n2002) );
  OAI221_X1 U972 ( .B1(n811), .B2(n1673), .C1(n779), .C2(n1674), .A(n2006), 
        .ZN(n2003) );
  NOR4_X1 U973 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .ZN(n1983) );
  OAI221_X1 U974 ( .B1(n42), .B2(n1683), .C1(n10), .C2(n1684), .A(n1991), .ZN(
        n1984) );
  OAI221_X1 U975 ( .B1(n938), .B2(n1678), .C1(n906), .C2(n1679), .A(n1990), 
        .ZN(n1985) );
  OAI221_X1 U976 ( .B1(n810), .B2(n1673), .C1(n778), .C2(n1674), .A(n1989), 
        .ZN(n1986) );
  NOR4_X1 U977 ( .A1(n1967), .A2(n1968), .A3(n1969), .A4(n1970), .ZN(n1966) );
  OAI221_X1 U978 ( .B1(n41), .B2(n1683), .C1(n9), .C2(n1684), .A(n1974), .ZN(
        n1967) );
  OAI221_X1 U979 ( .B1(n937), .B2(n1678), .C1(n905), .C2(n1679), .A(n1973), 
        .ZN(n1968) );
  OAI221_X1 U980 ( .B1(n809), .B2(n1673), .C1(n777), .C2(n1674), .A(n1972), 
        .ZN(n1969) );
  NOR4_X1 U981 ( .A1(n1950), .A2(n1951), .A3(n1952), .A4(n1953), .ZN(n1949) );
  OAI221_X1 U982 ( .B1(n40), .B2(n1683), .C1(n8), .C2(n1684), .A(n1957), .ZN(
        n1950) );
  OAI221_X1 U983 ( .B1(n936), .B2(n1678), .C1(n904), .C2(n1679), .A(n1956), 
        .ZN(n1951) );
  OAI221_X1 U984 ( .B1(n808), .B2(n1673), .C1(n776), .C2(n1674), .A(n1955), 
        .ZN(n1952) );
  NOR4_X1 U985 ( .A1(n1933), .A2(n1934), .A3(n1935), .A4(n1936), .ZN(n1932) );
  OAI221_X1 U986 ( .B1(n39), .B2(n1683), .C1(n7), .C2(n1684), .A(n1940), .ZN(
        n1933) );
  OAI221_X1 U987 ( .B1(n935), .B2(n1678), .C1(n903), .C2(n1679), .A(n1939), 
        .ZN(n1934) );
  OAI221_X1 U988 ( .B1(n807), .B2(n1673), .C1(n775), .C2(n1674), .A(n1938), 
        .ZN(n1935) );
  NOR4_X1 U989 ( .A1(n1916), .A2(n1917), .A3(n1918), .A4(n1919), .ZN(n1915) );
  OAI221_X1 U990 ( .B1(n38), .B2(n1683), .C1(n6), .C2(n1684), .A(n1923), .ZN(
        n1916) );
  OAI221_X1 U991 ( .B1(n934), .B2(n1678), .C1(n902), .C2(n1679), .A(n1922), 
        .ZN(n1917) );
  OAI221_X1 U992 ( .B1(n806), .B2(n1673), .C1(n774), .C2(n1674), .A(n1921), 
        .ZN(n1918) );
  NOR4_X1 U993 ( .A1(n1899), .A2(n1900), .A3(n1901), .A4(n1902), .ZN(n1898) );
  OAI221_X1 U994 ( .B1(n37), .B2(n1683), .C1(n5), .C2(n1684), .A(n1906), .ZN(
        n1899) );
  OAI221_X1 U995 ( .B1(n933), .B2(n1678), .C1(n901), .C2(n1679), .A(n1905), 
        .ZN(n1900) );
  OAI221_X1 U996 ( .B1(n805), .B2(n1673), .C1(n773), .C2(n1674), .A(n1904), 
        .ZN(n1901) );
  NOR4_X1 U997 ( .A1(n1882), .A2(n1883), .A3(n1884), .A4(n1885), .ZN(n1881) );
  OAI221_X1 U998 ( .B1(n36), .B2(n1683), .C1(n4), .C2(n1684), .A(n1889), .ZN(
        n1882) );
  OAI221_X1 U999 ( .B1(n932), .B2(n1678), .C1(n900), .C2(n1679), .A(n1888), 
        .ZN(n1883) );
  OAI221_X1 U1000 ( .B1(n804), .B2(n1673), .C1(n772), .C2(n1674), .A(n1887), 
        .ZN(n1884) );
  NOR4_X1 U1001 ( .A1(n1865), .A2(n1866), .A3(n1867), .A4(n1868), .ZN(n1864)
         );
  OAI221_X1 U1002 ( .B1(n35), .B2(n1683), .C1(n3), .C2(n1684), .A(n1872), .ZN(
        n1865) );
  OAI221_X1 U1003 ( .B1(n931), .B2(n1678), .C1(n899), .C2(n1679), .A(n1871), 
        .ZN(n1866) );
  OAI221_X1 U1004 ( .B1(n803), .B2(n1673), .C1(n771), .C2(n1674), .A(n1870), 
        .ZN(n1867) );
  NOR4_X1 U1005 ( .A1(n1831), .A2(n1832), .A3(n1833), .A4(n1834), .ZN(n1830)
         );
  OAI221_X1 U1006 ( .B1(n34), .B2(n1683), .C1(n2), .C2(n1684), .A(n1838), .ZN(
        n1831) );
  OAI221_X1 U1007 ( .B1(n930), .B2(n1678), .C1(n898), .C2(n1679), .A(n1837), 
        .ZN(n1832) );
  OAI221_X1 U1008 ( .B1(n802), .B2(n1673), .C1(n770), .C2(n1674), .A(n1836), 
        .ZN(n1833) );
  NOR4_X1 U1009 ( .A1(n1814), .A2(n1815), .A3(n1816), .A4(n1817), .ZN(n1813)
         );
  OAI221_X1 U1010 ( .B1(n33), .B2(n1683), .C1(n1), .C2(n1684), .A(n1821), .ZN(
        n1814) );
  OAI221_X1 U1011 ( .B1(n929), .B2(n1678), .C1(n897), .C2(n1679), .A(n1820), 
        .ZN(n1815) );
  OAI221_X1 U1012 ( .B1(n801), .B2(n1673), .C1(n769), .C2(n1674), .A(n1819), 
        .ZN(n1816) );
  NOR2_X1 U1013 ( .A1(n3715), .A2(wa[4]), .ZN(n2500) );
  INV_X1 U1014 ( .A(en_write), .ZN(n3715) );
  AOI22_X1 U1015 ( .A1(x23_s7_w[0]), .A2(n1086), .B1(x22_s6_w[0]), .B2(n1087), 
        .ZN(n1641) );
  AOI22_X1 U1016 ( .A1(x27_s11_w[0]), .A2(n1091), .B1(x26_s10_w[0]), .B2(n1092), .ZN(n1644) );
  AOI22_X1 U1017 ( .A1(x31_t6_w[0]), .A2(n1096), .B1(x30_t5_w[0]), .B2(n1097), 
        .ZN(n1647) );
  AOI22_X1 U1018 ( .A1(x23_s7_w[1]), .A2(n1086), .B1(x22_s6_w[1]), .B2(n1087), 
        .ZN(n1450) );
  AOI22_X1 U1019 ( .A1(x27_s11_w[1]), .A2(n1091), .B1(x26_s10_w[1]), .B2(n1092), .ZN(n1451) );
  AOI22_X1 U1020 ( .A1(x31_t6_w[1]), .A2(n1096), .B1(x30_t5_w[1]), .B2(n1097), 
        .ZN(n1452) );
  AOI22_X1 U1021 ( .A1(x23_s7_w[2]), .A2(n1086), .B1(x22_s6_w[2]), .B2(n1087), 
        .ZN(n1263) );
  AOI22_X1 U1022 ( .A1(x27_s11_w[2]), .A2(n1091), .B1(x26_s10_w[2]), .B2(n1092), .ZN(n1264) );
  AOI22_X1 U1023 ( .A1(x31_t6_w[2]), .A2(n1096), .B1(x30_t5_w[2]), .B2(n1097), 
        .ZN(n1265) );
  AOI22_X1 U1024 ( .A1(x23_s7_w[10]), .A2(n1086), .B1(x22_s6_w[10]), .B2(n1087), .ZN(n1620) );
  AOI22_X1 U1025 ( .A1(x27_s11_w[10]), .A2(n1091), .B1(x26_s10_w[10]), .B2(
        n1092), .ZN(n1621) );
  AOI22_X1 U1026 ( .A1(x31_t6_w[10]), .A2(n1096), .B1(x30_t5_w[10]), .B2(n1097), .ZN(n1622) );
  AOI22_X1 U1027 ( .A1(x23_s7_w[11]), .A2(n1086), .B1(x22_s6_w[11]), .B2(n1087), .ZN(n1603) );
  AOI22_X1 U1028 ( .A1(x27_s11_w[11]), .A2(n1091), .B1(x26_s10_w[11]), .B2(
        n1092), .ZN(n1604) );
  AOI22_X1 U1029 ( .A1(x31_t6_w[11]), .A2(n1096), .B1(x30_t5_w[11]), .B2(n1097), .ZN(n1605) );
  AOI22_X1 U1030 ( .A1(x23_s7_w[12]), .A2(n1086), .B1(x22_s6_w[12]), .B2(n1087), .ZN(n1586) );
  AOI22_X1 U1031 ( .A1(x27_s11_w[12]), .A2(n1091), .B1(x26_s10_w[12]), .B2(
        n1092), .ZN(n1587) );
  AOI22_X1 U1032 ( .A1(x31_t6_w[12]), .A2(n1096), .B1(x30_t5_w[12]), .B2(n1097), .ZN(n1588) );
  AOI22_X1 U1033 ( .A1(x23_s7_w[13]), .A2(n1086), .B1(x22_s6_w[13]), .B2(n1087), .ZN(n1569) );
  AOI22_X1 U1034 ( .A1(x27_s11_w[13]), .A2(n1091), .B1(x26_s10_w[13]), .B2(
        n1092), .ZN(n1570) );
  AOI22_X1 U1035 ( .A1(x31_t6_w[13]), .A2(n1096), .B1(x30_t5_w[13]), .B2(n1097), .ZN(n1571) );
  AOI22_X1 U1036 ( .A1(x23_s7_w[14]), .A2(n1086), .B1(x22_s6_w[14]), .B2(n1087), .ZN(n1552) );
  AOI22_X1 U1037 ( .A1(x27_s11_w[14]), .A2(n1091), .B1(x26_s10_w[14]), .B2(
        n1092), .ZN(n1553) );
  AOI22_X1 U1038 ( .A1(x31_t6_w[14]), .A2(n1096), .B1(x30_t5_w[14]), .B2(n1097), .ZN(n1554) );
  AOI22_X1 U1039 ( .A1(x23_s7_w[15]), .A2(n1086), .B1(x22_s6_w[15]), .B2(n1087), .ZN(n1535) );
  AOI22_X1 U1040 ( .A1(x27_s11_w[15]), .A2(n1091), .B1(x26_s10_w[15]), .B2(
        n1092), .ZN(n1536) );
  AOI22_X1 U1041 ( .A1(x31_t6_w[15]), .A2(n1096), .B1(x30_t5_w[15]), .B2(n1097), .ZN(n1537) );
  AOI22_X1 U1042 ( .A1(x23_s7_w[16]), .A2(n1086), .B1(x22_s6_w[16]), .B2(n1087), .ZN(n1518) );
  AOI22_X1 U1043 ( .A1(x27_s11_w[16]), .A2(n1091), .B1(x26_s10_w[16]), .B2(
        n1092), .ZN(n1519) );
  AOI22_X1 U1044 ( .A1(x31_t6_w[16]), .A2(n1096), .B1(x30_t5_w[16]), .B2(n1097), .ZN(n1520) );
  AOI22_X1 U1045 ( .A1(x23_s7_w[17]), .A2(n1086), .B1(x22_s6_w[17]), .B2(n1087), .ZN(n1501) );
  AOI22_X1 U1046 ( .A1(x27_s11_w[17]), .A2(n1091), .B1(x26_s10_w[17]), .B2(
        n1092), .ZN(n1502) );
  AOI22_X1 U1047 ( .A1(x31_t6_w[17]), .A2(n1096), .B1(x30_t5_w[17]), .B2(n1097), .ZN(n1503) );
  AOI22_X1 U1048 ( .A1(x23_s7_w[18]), .A2(n1086), .B1(x22_s6_w[18]), .B2(n1087), .ZN(n1484) );
  AOI22_X1 U1049 ( .A1(x27_s11_w[18]), .A2(n1091), .B1(x26_s10_w[18]), .B2(
        n1092), .ZN(n1485) );
  AOI22_X1 U1050 ( .A1(x31_t6_w[18]), .A2(n1096), .B1(x30_t5_w[18]), .B2(n1097), .ZN(n1486) );
  AOI22_X1 U1051 ( .A1(x23_s7_w[19]), .A2(n1086), .B1(x22_s6_w[19]), .B2(n1087), .ZN(n1467) );
  AOI22_X1 U1052 ( .A1(x27_s11_w[19]), .A2(n1091), .B1(x26_s10_w[19]), .B2(
        n1092), .ZN(n1468) );
  AOI22_X1 U1053 ( .A1(x31_t6_w[19]), .A2(n1096), .B1(x30_t5_w[19]), .B2(n1097), .ZN(n1469) );
  AOI22_X1 U1054 ( .A1(x23_s7_w[20]), .A2(n1086), .B1(x22_s6_w[20]), .B2(n1087), .ZN(n1433) );
  AOI22_X1 U1055 ( .A1(x27_s11_w[20]), .A2(n1091), .B1(x26_s10_w[20]), .B2(
        n1092), .ZN(n1434) );
  AOI22_X1 U1056 ( .A1(x31_t6_w[20]), .A2(n1096), .B1(x30_t5_w[20]), .B2(n1097), .ZN(n1435) );
  AOI22_X1 U1057 ( .A1(x23_s7_w[21]), .A2(n1086), .B1(x22_s6_w[21]), .B2(n1087), .ZN(n1416) );
  AOI22_X1 U1058 ( .A1(x27_s11_w[21]), .A2(n1091), .B1(x26_s10_w[21]), .B2(
        n1092), .ZN(n1417) );
  AOI22_X1 U1059 ( .A1(x31_t6_w[21]), .A2(n1096), .B1(x30_t5_w[21]), .B2(n1097), .ZN(n1418) );
  AOI22_X1 U1060 ( .A1(x23_s7_w[22]), .A2(n1086), .B1(x22_s6_w[22]), .B2(n1087), .ZN(n1399) );
  AOI22_X1 U1061 ( .A1(x27_s11_w[22]), .A2(n1091), .B1(x26_s10_w[22]), .B2(
        n1092), .ZN(n1400) );
  AOI22_X1 U1062 ( .A1(x31_t6_w[22]), .A2(n1096), .B1(x30_t5_w[22]), .B2(n1097), .ZN(n1401) );
  AOI22_X1 U1063 ( .A1(x23_s7_w[23]), .A2(n1086), .B1(x22_s6_w[23]), .B2(n1087), .ZN(n1382) );
  AOI22_X1 U1064 ( .A1(x27_s11_w[23]), .A2(n1091), .B1(x26_s10_w[23]), .B2(
        n1092), .ZN(n1383) );
  AOI22_X1 U1065 ( .A1(x31_t6_w[23]), .A2(n1096), .B1(x30_t5_w[23]), .B2(n1097), .ZN(n1384) );
  AOI22_X1 U1066 ( .A1(x23_s7_w[24]), .A2(n1086), .B1(x22_s6_w[24]), .B2(n1087), .ZN(n1365) );
  AOI22_X1 U1067 ( .A1(x27_s11_w[24]), .A2(n1091), .B1(x26_s10_w[24]), .B2(
        n1092), .ZN(n1366) );
  AOI22_X1 U1068 ( .A1(x31_t6_w[24]), .A2(n1096), .B1(x30_t5_w[24]), .B2(n1097), .ZN(n1367) );
  AOI22_X1 U1069 ( .A1(x23_s7_w[25]), .A2(n1086), .B1(x22_s6_w[25]), .B2(n1087), .ZN(n1348) );
  AOI22_X1 U1070 ( .A1(x27_s11_w[25]), .A2(n1091), .B1(x26_s10_w[25]), .B2(
        n1092), .ZN(n1349) );
  AOI22_X1 U1071 ( .A1(x31_t6_w[25]), .A2(n1096), .B1(x30_t5_w[25]), .B2(n1097), .ZN(n1350) );
  AOI22_X1 U1072 ( .A1(x23_s7_w[26]), .A2(n1086), .B1(x22_s6_w[26]), .B2(n1087), .ZN(n1331) );
  AOI22_X1 U1073 ( .A1(x27_s11_w[26]), .A2(n1091), .B1(x26_s10_w[26]), .B2(
        n1092), .ZN(n1332) );
  AOI22_X1 U1074 ( .A1(x31_t6_w[26]), .A2(n1096), .B1(x30_t5_w[26]), .B2(n1097), .ZN(n1333) );
  AOI22_X1 U1075 ( .A1(x23_s7_w[27]), .A2(n1086), .B1(x22_s6_w[27]), .B2(n1087), .ZN(n1314) );
  AOI22_X1 U1076 ( .A1(x27_s11_w[27]), .A2(n1091), .B1(x26_s10_w[27]), .B2(
        n1092), .ZN(n1315) );
  AOI22_X1 U1077 ( .A1(x31_t6_w[27]), .A2(n1096), .B1(x30_t5_w[27]), .B2(n1097), .ZN(n1316) );
  AOI22_X1 U1078 ( .A1(x23_s7_w[28]), .A2(n1086), .B1(x22_s6_w[28]), .B2(n1087), .ZN(n1297) );
  AOI22_X1 U1079 ( .A1(x27_s11_w[28]), .A2(n1091), .B1(x26_s10_w[28]), .B2(
        n1092), .ZN(n1298) );
  AOI22_X1 U1080 ( .A1(x31_t6_w[28]), .A2(n1096), .B1(x30_t5_w[28]), .B2(n1097), .ZN(n1299) );
  AOI22_X1 U1081 ( .A1(x23_s7_w[29]), .A2(n1086), .B1(x22_s6_w[29]), .B2(n1087), .ZN(n1280) );
  AOI22_X1 U1082 ( .A1(x27_s11_w[29]), .A2(n1091), .B1(x26_s10_w[29]), .B2(
        n1092), .ZN(n1281) );
  AOI22_X1 U1083 ( .A1(x31_t6_w[29]), .A2(n1096), .B1(x30_t5_w[29]), .B2(n1097), .ZN(n1282) );
  AOI22_X1 U1084 ( .A1(x23_s7_w[30]), .A2(n1086), .B1(x22_s6_w[30]), .B2(n1087), .ZN(n1246) );
  AOI22_X1 U1085 ( .A1(x27_s11_w[30]), .A2(n1091), .B1(x26_s10_w[30]), .B2(
        n1092), .ZN(n1247) );
  AOI22_X1 U1086 ( .A1(x31_t6_w[30]), .A2(n1096), .B1(x30_t5_w[30]), .B2(n1097), .ZN(n1248) );
  AOI22_X1 U1087 ( .A1(x23_s7_w[3]), .A2(n1086), .B1(x22_s6_w[3]), .B2(n1087), 
        .ZN(n1212) );
  AOI22_X1 U1088 ( .A1(x27_s11_w[3]), .A2(n1091), .B1(x26_s10_w[3]), .B2(n1092), .ZN(n1213) );
  AOI22_X1 U1089 ( .A1(x31_t6_w[3]), .A2(n1096), .B1(x30_t5_w[3]), .B2(n1097), 
        .ZN(n1214) );
  AOI22_X1 U1090 ( .A1(x23_s7_w[4]), .A2(n1086), .B1(x22_s6_w[4]), .B2(n1087), 
        .ZN(n1195) );
  AOI22_X1 U1091 ( .A1(x27_s11_w[4]), .A2(n1091), .B1(x26_s10_w[4]), .B2(n1092), .ZN(n1196) );
  AOI22_X1 U1092 ( .A1(x31_t6_w[4]), .A2(n1096), .B1(x30_t5_w[4]), .B2(n1097), 
        .ZN(n1197) );
  AOI22_X1 U1093 ( .A1(x23_s7_w[5]), .A2(n1086), .B1(x22_s6_w[5]), .B2(n1087), 
        .ZN(n1178) );
  AOI22_X1 U1094 ( .A1(x27_s11_w[5]), .A2(n1091), .B1(x26_s10_w[5]), .B2(n1092), .ZN(n1179) );
  AOI22_X1 U1095 ( .A1(x31_t6_w[5]), .A2(n1096), .B1(x30_t5_w[5]), .B2(n1097), 
        .ZN(n1180) );
  AOI22_X1 U1096 ( .A1(x23_s7_w[6]), .A2(n1086), .B1(x22_s6_w[6]), .B2(n1087), 
        .ZN(n1161) );
  AOI22_X1 U1097 ( .A1(x27_s11_w[6]), .A2(n1091), .B1(x26_s10_w[6]), .B2(n1092), .ZN(n1162) );
  AOI22_X1 U1098 ( .A1(x31_t6_w[6]), .A2(n1096), .B1(x30_t5_w[6]), .B2(n1097), 
        .ZN(n1163) );
  AOI22_X1 U1099 ( .A1(x23_s7_w[7]), .A2(n1086), .B1(x22_s6_w[7]), .B2(n1087), 
        .ZN(n1144) );
  AOI22_X1 U1100 ( .A1(x27_s11_w[7]), .A2(n1091), .B1(x26_s10_w[7]), .B2(n1092), .ZN(n1145) );
  AOI22_X1 U1101 ( .A1(x31_t6_w[7]), .A2(n1096), .B1(x30_t5_w[7]), .B2(n1097), 
        .ZN(n1146) );
  AOI22_X1 U1102 ( .A1(x23_s7_w[8]), .A2(n1086), .B1(x22_s6_w[8]), .B2(n1087), 
        .ZN(n1127) );
  AOI22_X1 U1103 ( .A1(x27_s11_w[8]), .A2(n1091), .B1(x26_s10_w[8]), .B2(n1092), .ZN(n1128) );
  AOI22_X1 U1104 ( .A1(x31_t6_w[8]), .A2(n1096), .B1(x30_t5_w[8]), .B2(n1097), 
        .ZN(n1129) );
  AOI22_X1 U1105 ( .A1(x23_s7_w[9]), .A2(n1086), .B1(x22_s6_w[9]), .B2(n1087), 
        .ZN(n1085) );
  AOI22_X1 U1106 ( .A1(x27_s11_w[9]), .A2(n1091), .B1(x26_s10_w[9]), .B2(n1092), .ZN(n1090) );
  AOI22_X1 U1107 ( .A1(x31_t6_w[9]), .A2(n1096), .B1(x30_t5_w[9]), .B2(n1097), 
        .ZN(n1095) );
  AOI22_X1 U1108 ( .A1(x23_s7_w[31]), .A2(n1086), .B1(x22_s6_w[31]), .B2(n1087), .ZN(n1229) );
  AOI22_X1 U1109 ( .A1(x27_s11_w[31]), .A2(n1091), .B1(x26_s10_w[31]), .B2(
        n1092), .ZN(n1230) );
  AOI22_X1 U1110 ( .A1(x31_t6_w[31]), .A2(n1096), .B1(x30_t5_w[31]), .B2(n1097), .ZN(n1231) );
  AOI22_X1 U1111 ( .A1(n1676), .A2(x23_s7_w[0]), .B1(n1677), .B2(x22_s6_w[0]), 
        .ZN(n2231) );
  AOI22_X1 U1112 ( .A1(n1681), .A2(x27_s11_w[0]), .B1(n1682), .B2(x26_s10_w[0]), .ZN(n2234) );
  AOI22_X1 U1113 ( .A1(n1686), .A2(x31_t6_w[0]), .B1(n1687), .B2(x30_t5_w[0]), 
        .ZN(n2237) );
  AOI22_X1 U1114 ( .A1(n1676), .A2(x23_s7_w[1]), .B1(n1677), .B2(x22_s6_w[1]), 
        .ZN(n2040) );
  AOI22_X1 U1115 ( .A1(n1681), .A2(x27_s11_w[1]), .B1(n1682), .B2(x26_s10_w[1]), .ZN(n2041) );
  AOI22_X1 U1116 ( .A1(n1686), .A2(x31_t6_w[1]), .B1(n1687), .B2(x30_t5_w[1]), 
        .ZN(n2042) );
  AOI22_X1 U1117 ( .A1(n1676), .A2(x23_s7_w[2]), .B1(n1677), .B2(x22_s6_w[2]), 
        .ZN(n1853) );
  AOI22_X1 U1118 ( .A1(n1681), .A2(x27_s11_w[2]), .B1(n1682), .B2(x26_s10_w[2]), .ZN(n1854) );
  AOI22_X1 U1119 ( .A1(n1686), .A2(x31_t6_w[2]), .B1(n1687), .B2(x30_t5_w[2]), 
        .ZN(n1855) );
  AOI22_X1 U1120 ( .A1(n1676), .A2(x23_s7_w[3]), .B1(n1677), .B2(x22_s6_w[3]), 
        .ZN(n1802) );
  AOI22_X1 U1121 ( .A1(n1681), .A2(x27_s11_w[3]), .B1(n1682), .B2(x26_s10_w[3]), .ZN(n1803) );
  AOI22_X1 U1122 ( .A1(n1686), .A2(x31_t6_w[3]), .B1(n1687), .B2(x30_t5_w[3]), 
        .ZN(n1804) );
  AOI22_X1 U1123 ( .A1(n1676), .A2(x23_s7_w[4]), .B1(n1677), .B2(x22_s6_w[4]), 
        .ZN(n1785) );
  AOI22_X1 U1124 ( .A1(n1681), .A2(x27_s11_w[4]), .B1(n1682), .B2(x26_s10_w[4]), .ZN(n1786) );
  AOI22_X1 U1125 ( .A1(n1686), .A2(x31_t6_w[4]), .B1(n1687), .B2(x30_t5_w[4]), 
        .ZN(n1787) );
  AOI22_X1 U1126 ( .A1(n1676), .A2(x23_s7_w[5]), .B1(n1677), .B2(x22_s6_w[5]), 
        .ZN(n1768) );
  AOI22_X1 U1127 ( .A1(n1681), .A2(x27_s11_w[5]), .B1(n1682), .B2(x26_s10_w[5]), .ZN(n1769) );
  AOI22_X1 U1128 ( .A1(n1686), .A2(x31_t6_w[5]), .B1(n1687), .B2(x30_t5_w[5]), 
        .ZN(n1770) );
  AOI22_X1 U1129 ( .A1(n1676), .A2(x23_s7_w[6]), .B1(n1677), .B2(x22_s6_w[6]), 
        .ZN(n1751) );
  AOI22_X1 U1130 ( .A1(n1681), .A2(x27_s11_w[6]), .B1(n1682), .B2(x26_s10_w[6]), .ZN(n1752) );
  AOI22_X1 U1131 ( .A1(n1686), .A2(x31_t6_w[6]), .B1(n1687), .B2(x30_t5_w[6]), 
        .ZN(n1753) );
  AOI22_X1 U1132 ( .A1(n1676), .A2(x23_s7_w[7]), .B1(n1677), .B2(x22_s6_w[7]), 
        .ZN(n1734) );
  AOI22_X1 U1133 ( .A1(n1681), .A2(x27_s11_w[7]), .B1(n1682), .B2(x26_s10_w[7]), .ZN(n1735) );
  AOI22_X1 U1134 ( .A1(n1686), .A2(x31_t6_w[7]), .B1(n1687), .B2(x30_t5_w[7]), 
        .ZN(n1736) );
  AOI22_X1 U1135 ( .A1(n1676), .A2(x23_s7_w[8]), .B1(n1677), .B2(x22_s6_w[8]), 
        .ZN(n1717) );
  AOI22_X1 U1136 ( .A1(n1681), .A2(x27_s11_w[8]), .B1(n1682), .B2(x26_s10_w[8]), .ZN(n1718) );
  AOI22_X1 U1137 ( .A1(n1686), .A2(x31_t6_w[8]), .B1(n1687), .B2(x30_t5_w[8]), 
        .ZN(n1719) );
  AOI22_X1 U1138 ( .A1(n1676), .A2(x23_s7_w[9]), .B1(n1677), .B2(x22_s6_w[9]), 
        .ZN(n1675) );
  AOI22_X1 U1139 ( .A1(n1681), .A2(x27_s11_w[9]), .B1(n1682), .B2(x26_s10_w[9]), .ZN(n1680) );
  AOI22_X1 U1140 ( .A1(n1686), .A2(x31_t6_w[9]), .B1(n1687), .B2(x30_t5_w[9]), 
        .ZN(n1685) );
  AOI22_X1 U1141 ( .A1(n1676), .A2(x23_s7_w[10]), .B1(n1677), .B2(x22_s6_w[10]), .ZN(n2210) );
  AOI22_X1 U1142 ( .A1(n1681), .A2(x27_s11_w[10]), .B1(n1682), .B2(
        x26_s10_w[10]), .ZN(n2211) );
  AOI22_X1 U1143 ( .A1(n1686), .A2(x31_t6_w[10]), .B1(n1687), .B2(x30_t5_w[10]), .ZN(n2212) );
  AOI22_X1 U1144 ( .A1(n1676), .A2(x23_s7_w[11]), .B1(n1677), .B2(x22_s6_w[11]), .ZN(n2193) );
  AOI22_X1 U1145 ( .A1(n1681), .A2(x27_s11_w[11]), .B1(n1682), .B2(
        x26_s10_w[11]), .ZN(n2194) );
  AOI22_X1 U1146 ( .A1(n1686), .A2(x31_t6_w[11]), .B1(n1687), .B2(x30_t5_w[11]), .ZN(n2195) );
  AOI22_X1 U1147 ( .A1(n1676), .A2(x23_s7_w[12]), .B1(n1677), .B2(x22_s6_w[12]), .ZN(n2176) );
  AOI22_X1 U1148 ( .A1(n1681), .A2(x27_s11_w[12]), .B1(n1682), .B2(
        x26_s10_w[12]), .ZN(n2177) );
  AOI22_X1 U1149 ( .A1(n1686), .A2(x31_t6_w[12]), .B1(n1687), .B2(x30_t5_w[12]), .ZN(n2178) );
  AOI22_X1 U1150 ( .A1(n1676), .A2(x23_s7_w[13]), .B1(n1677), .B2(x22_s6_w[13]), .ZN(n2159) );
  AOI22_X1 U1151 ( .A1(n1681), .A2(x27_s11_w[13]), .B1(n1682), .B2(
        x26_s10_w[13]), .ZN(n2160) );
  AOI22_X1 U1152 ( .A1(n1686), .A2(x31_t6_w[13]), .B1(n1687), .B2(x30_t5_w[13]), .ZN(n2161) );
  AOI22_X1 U1153 ( .A1(n1676), .A2(x23_s7_w[14]), .B1(n1677), .B2(x22_s6_w[14]), .ZN(n2142) );
  AOI22_X1 U1154 ( .A1(n1681), .A2(x27_s11_w[14]), .B1(n1682), .B2(
        x26_s10_w[14]), .ZN(n2143) );
  AOI22_X1 U1155 ( .A1(n1686), .A2(x31_t6_w[14]), .B1(n1687), .B2(x30_t5_w[14]), .ZN(n2144) );
  AOI22_X1 U1156 ( .A1(n1676), .A2(x23_s7_w[15]), .B1(n1677), .B2(x22_s6_w[15]), .ZN(n2125) );
  AOI22_X1 U1157 ( .A1(n1681), .A2(x27_s11_w[15]), .B1(n1682), .B2(
        x26_s10_w[15]), .ZN(n2126) );
  AOI22_X1 U1158 ( .A1(n1686), .A2(x31_t6_w[15]), .B1(n1687), .B2(x30_t5_w[15]), .ZN(n2127) );
  AOI22_X1 U1159 ( .A1(n1676), .A2(x23_s7_w[16]), .B1(n1677), .B2(x22_s6_w[16]), .ZN(n2108) );
  AOI22_X1 U1160 ( .A1(n1681), .A2(x27_s11_w[16]), .B1(n1682), .B2(
        x26_s10_w[16]), .ZN(n2109) );
  AOI22_X1 U1161 ( .A1(n1686), .A2(x31_t6_w[16]), .B1(n1687), .B2(x30_t5_w[16]), .ZN(n2110) );
  AOI22_X1 U1162 ( .A1(n1676), .A2(x23_s7_w[17]), .B1(n1677), .B2(x22_s6_w[17]), .ZN(n2091) );
  AOI22_X1 U1163 ( .A1(n1681), .A2(x27_s11_w[17]), .B1(n1682), .B2(
        x26_s10_w[17]), .ZN(n2092) );
  AOI22_X1 U1164 ( .A1(n1686), .A2(x31_t6_w[17]), .B1(n1687), .B2(x30_t5_w[17]), .ZN(n2093) );
  AOI22_X1 U1165 ( .A1(n1676), .A2(x23_s7_w[18]), .B1(n1677), .B2(x22_s6_w[18]), .ZN(n2074) );
  AOI22_X1 U1166 ( .A1(n1681), .A2(x27_s11_w[18]), .B1(n1682), .B2(
        x26_s10_w[18]), .ZN(n2075) );
  AOI22_X1 U1167 ( .A1(n1686), .A2(x31_t6_w[18]), .B1(n1687), .B2(x30_t5_w[18]), .ZN(n2076) );
  AOI22_X1 U1168 ( .A1(n1676), .A2(x23_s7_w[19]), .B1(n1677), .B2(x22_s6_w[19]), .ZN(n2057) );
  AOI22_X1 U1169 ( .A1(n1681), .A2(x27_s11_w[19]), .B1(n1682), .B2(
        x26_s10_w[19]), .ZN(n2058) );
  AOI22_X1 U1170 ( .A1(n1686), .A2(x31_t6_w[19]), .B1(n1687), .B2(x30_t5_w[19]), .ZN(n2059) );
  AOI22_X1 U1171 ( .A1(n1676), .A2(x23_s7_w[20]), .B1(n1677), .B2(x22_s6_w[20]), .ZN(n2023) );
  AOI22_X1 U1172 ( .A1(n1681), .A2(x27_s11_w[20]), .B1(n1682), .B2(
        x26_s10_w[20]), .ZN(n2024) );
  AOI22_X1 U1173 ( .A1(n1686), .A2(x31_t6_w[20]), .B1(n1687), .B2(x30_t5_w[20]), .ZN(n2025) );
  AOI22_X1 U1174 ( .A1(n1676), .A2(x23_s7_w[21]), .B1(n1677), .B2(x22_s6_w[21]), .ZN(n2006) );
  AOI22_X1 U1175 ( .A1(n1681), .A2(x27_s11_w[21]), .B1(n1682), .B2(
        x26_s10_w[21]), .ZN(n2007) );
  AOI22_X1 U1176 ( .A1(n1686), .A2(x31_t6_w[21]), .B1(n1687), .B2(x30_t5_w[21]), .ZN(n2008) );
  AOI22_X1 U1177 ( .A1(n1676), .A2(x23_s7_w[22]), .B1(n1677), .B2(x22_s6_w[22]), .ZN(n1989) );
  AOI22_X1 U1178 ( .A1(n1681), .A2(x27_s11_w[22]), .B1(n1682), .B2(
        x26_s10_w[22]), .ZN(n1990) );
  AOI22_X1 U1179 ( .A1(n1686), .A2(x31_t6_w[22]), .B1(n1687), .B2(x30_t5_w[22]), .ZN(n1991) );
  AOI22_X1 U1180 ( .A1(n1676), .A2(x23_s7_w[23]), .B1(n1677), .B2(x22_s6_w[23]), .ZN(n1972) );
  AOI22_X1 U1181 ( .A1(n1681), .A2(x27_s11_w[23]), .B1(n1682), .B2(
        x26_s10_w[23]), .ZN(n1973) );
  AOI22_X1 U1182 ( .A1(n1686), .A2(x31_t6_w[23]), .B1(n1687), .B2(x30_t5_w[23]), .ZN(n1974) );
  AOI22_X1 U1183 ( .A1(n1676), .A2(x23_s7_w[24]), .B1(n1677), .B2(x22_s6_w[24]), .ZN(n1955) );
  AOI22_X1 U1184 ( .A1(n1681), .A2(x27_s11_w[24]), .B1(n1682), .B2(
        x26_s10_w[24]), .ZN(n1956) );
  AOI22_X1 U1185 ( .A1(n1686), .A2(x31_t6_w[24]), .B1(n1687), .B2(x30_t5_w[24]), .ZN(n1957) );
  AOI22_X1 U1186 ( .A1(n1676), .A2(x23_s7_w[25]), .B1(n1677), .B2(x22_s6_w[25]), .ZN(n1938) );
  AOI22_X1 U1187 ( .A1(n1681), .A2(x27_s11_w[25]), .B1(n1682), .B2(
        x26_s10_w[25]), .ZN(n1939) );
  AOI22_X1 U1188 ( .A1(n1686), .A2(x31_t6_w[25]), .B1(n1687), .B2(x30_t5_w[25]), .ZN(n1940) );
  AOI22_X1 U1189 ( .A1(n1676), .A2(x23_s7_w[26]), .B1(n1677), .B2(x22_s6_w[26]), .ZN(n1921) );
  AOI22_X1 U1190 ( .A1(n1681), .A2(x27_s11_w[26]), .B1(n1682), .B2(
        x26_s10_w[26]), .ZN(n1922) );
  AOI22_X1 U1191 ( .A1(n1686), .A2(x31_t6_w[26]), .B1(n1687), .B2(x30_t5_w[26]), .ZN(n1923) );
  AOI22_X1 U1192 ( .A1(n1676), .A2(x23_s7_w[27]), .B1(n1677), .B2(x22_s6_w[27]), .ZN(n1904) );
  AOI22_X1 U1193 ( .A1(n1681), .A2(x27_s11_w[27]), .B1(n1682), .B2(
        x26_s10_w[27]), .ZN(n1905) );
  AOI22_X1 U1194 ( .A1(n1686), .A2(x31_t6_w[27]), .B1(n1687), .B2(x30_t5_w[27]), .ZN(n1906) );
  AOI22_X1 U1195 ( .A1(n1676), .A2(x23_s7_w[28]), .B1(n1677), .B2(x22_s6_w[28]), .ZN(n1887) );
  AOI22_X1 U1196 ( .A1(n1681), .A2(x27_s11_w[28]), .B1(n1682), .B2(
        x26_s10_w[28]), .ZN(n1888) );
  AOI22_X1 U1197 ( .A1(n1686), .A2(x31_t6_w[28]), .B1(n1687), .B2(x30_t5_w[28]), .ZN(n1889) );
  AOI22_X1 U1198 ( .A1(n1676), .A2(x23_s7_w[29]), .B1(n1677), .B2(x22_s6_w[29]), .ZN(n1870) );
  AOI22_X1 U1199 ( .A1(n1681), .A2(x27_s11_w[29]), .B1(n1682), .B2(
        x26_s10_w[29]), .ZN(n1871) );
  AOI22_X1 U1200 ( .A1(n1686), .A2(x31_t6_w[29]), .B1(n1687), .B2(x30_t5_w[29]), .ZN(n1872) );
  AOI22_X1 U1201 ( .A1(n1676), .A2(x23_s7_w[30]), .B1(n1677), .B2(x22_s6_w[30]), .ZN(n1836) );
  AOI22_X1 U1202 ( .A1(n1681), .A2(x27_s11_w[30]), .B1(n1682), .B2(
        x26_s10_w[30]), .ZN(n1837) );
  AOI22_X1 U1203 ( .A1(n1686), .A2(x31_t6_w[30]), .B1(n1687), .B2(x30_t5_w[30]), .ZN(n1838) );
  AOI22_X1 U1204 ( .A1(n1676), .A2(x23_s7_w[31]), .B1(n1677), .B2(x22_s6_w[31]), .ZN(n1819) );
  AOI22_X1 U1205 ( .A1(n1681), .A2(x27_s11_w[31]), .B1(n1682), .B2(
        x26_s10_w[31]), .ZN(n1820) );
  AOI22_X1 U1206 ( .A1(n1686), .A2(x31_t6_w[31]), .B1(n1687), .B2(x30_t5_w[31]), .ZN(n1821) );
  OAI221_X1 U1207 ( .B1(n1078), .B2(n765), .C1(n1079), .C2(n733), .A(n1211), 
        .ZN(n1210) );
  AOI22_X1 U1208 ( .A1(x17_a7_w[3]), .A2(n1081), .B1(x16_a6_w[3]), .B2(n1082), 
        .ZN(n1211) );
  OAI221_X1 U1209 ( .B1(n1103), .B2(n317), .C1(n1104), .C2(n285), .A(n1217), 
        .ZN(n1215) );
  AOI22_X1 U1210 ( .A1(x7_t2_w[3]), .A2(n1106), .B1(x6_t1_w[3]), .B2(n1107), 
        .ZN(n1217) );
  OAI221_X1 U1211 ( .B1(n1078), .B2(n764), .C1(n1079), .C2(n732), .A(n1194), 
        .ZN(n1193) );
  AOI22_X1 U1212 ( .A1(x17_a7_w[4]), .A2(n1081), .B1(x16_a6_w[4]), .B2(n1082), 
        .ZN(n1194) );
  OAI221_X1 U1213 ( .B1(n1103), .B2(n316), .C1(n1104), .C2(n284), .A(n1200), 
        .ZN(n1198) );
  AOI22_X1 U1214 ( .A1(x7_t2_w[4]), .A2(n1106), .B1(x6_t1_w[4]), .B2(n1107), 
        .ZN(n1200) );
  OAI221_X1 U1215 ( .B1(n1078), .B2(n763), .C1(n1079), .C2(n731), .A(n1177), 
        .ZN(n1176) );
  AOI22_X1 U1216 ( .A1(x17_a7_w[5]), .A2(n1081), .B1(x16_a6_w[5]), .B2(n1082), 
        .ZN(n1177) );
  OAI221_X1 U1217 ( .B1(n1103), .B2(n315), .C1(n1104), .C2(n283), .A(n1183), 
        .ZN(n1181) );
  AOI22_X1 U1218 ( .A1(x7_t2_w[5]), .A2(n1106), .B1(x6_t1_w[5]), .B2(n1107), 
        .ZN(n1183) );
  OAI221_X1 U1219 ( .B1(n1078), .B2(n762), .C1(n1079), .C2(n730), .A(n1160), 
        .ZN(n1159) );
  AOI22_X1 U1220 ( .A1(x17_a7_w[6]), .A2(n1081), .B1(x16_a6_w[6]), .B2(n1082), 
        .ZN(n1160) );
  OAI221_X1 U1221 ( .B1(n1103), .B2(n314), .C1(n1104), .C2(n282), .A(n1166), 
        .ZN(n1164) );
  AOI22_X1 U1222 ( .A1(x7_t2_w[6]), .A2(n1106), .B1(x6_t1_w[6]), .B2(n1107), 
        .ZN(n1166) );
  OAI221_X1 U1223 ( .B1(n1078), .B2(n761), .C1(n1079), .C2(n729), .A(n1143), 
        .ZN(n1142) );
  AOI22_X1 U1224 ( .A1(x17_a7_w[7]), .A2(n1081), .B1(x16_a6_w[7]), .B2(n1082), 
        .ZN(n1143) );
  OAI221_X1 U1225 ( .B1(n1103), .B2(n313), .C1(n1104), .C2(n281), .A(n1149), 
        .ZN(n1147) );
  AOI22_X1 U1226 ( .A1(x7_t2_w[7]), .A2(n1106), .B1(x6_t1_w[7]), .B2(n1107), 
        .ZN(n1149) );
  OAI221_X1 U1227 ( .B1(n1078), .B2(n760), .C1(n1079), .C2(n728), .A(n1126), 
        .ZN(n1125) );
  AOI22_X1 U1228 ( .A1(x17_a7_w[8]), .A2(n1081), .B1(x16_a6_w[8]), .B2(n1082), 
        .ZN(n1126) );
  OAI221_X1 U1229 ( .B1(n1103), .B2(n312), .C1(n1104), .C2(n280), .A(n1132), 
        .ZN(n1130) );
  AOI22_X1 U1230 ( .A1(x7_t2_w[8]), .A2(n1106), .B1(x6_t1_w[8]), .B2(n1107), 
        .ZN(n1132) );
  OAI221_X1 U1231 ( .B1(n1078), .B2(n759), .C1(n1079), .C2(n727), .A(n1080), 
        .ZN(n1077) );
  AOI22_X1 U1232 ( .A1(x17_a7_w[9]), .A2(n1081), .B1(x16_a6_w[9]), .B2(n1082), 
        .ZN(n1080) );
  OAI221_X1 U1233 ( .B1(n1103), .B2(n311), .C1(n1104), .C2(n279), .A(n1105), 
        .ZN(n1099) );
  AOI22_X1 U1234 ( .A1(x7_t2_w[9]), .A2(n1106), .B1(x6_t1_w[9]), .B2(n1107), 
        .ZN(n1105) );
  OAI221_X1 U1235 ( .B1(n1078), .B2(n737), .C1(n1079), .C2(n705), .A(n1228), 
        .ZN(n1227) );
  AOI22_X1 U1236 ( .A1(x17_a7_w[31]), .A2(n1081), .B1(x16_a6_w[31]), .B2(n1082), .ZN(n1228) );
  OAI221_X1 U1237 ( .B1(n1103), .B2(n289), .C1(n1104), .C2(n257), .A(n1234), 
        .ZN(n1232) );
  AOI22_X1 U1238 ( .A1(x7_t2_w[31]), .A2(n1106), .B1(x6_t1_w[31]), .B2(n1107), 
        .ZN(n1234) );
  OAI221_X1 U1239 ( .B1(n768), .B2(n1668), .C1(n736), .C2(n1669), .A(n2226), 
        .ZN(n2225) );
  AOI22_X1 U1240 ( .A1(n1671), .A2(x17_a7_w[0]), .B1(n1672), .B2(x16_a6_w[0]), 
        .ZN(n2226) );
  OAI221_X1 U1241 ( .B1(n320), .B2(n1693), .C1(n288), .C2(n1694), .A(n2245), 
        .ZN(n2240) );
  AOI22_X1 U1242 ( .A1(n1696), .A2(x7_t2_w[0]), .B1(n1697), .B2(x6_t1_w[0]), 
        .ZN(n2245) );
  OAI221_X1 U1243 ( .B1(n767), .B2(n1668), .C1(n735), .C2(n1669), .A(n2039), 
        .ZN(n2038) );
  AOI22_X1 U1244 ( .A1(n1671), .A2(x17_a7_w[1]), .B1(n1672), .B2(x16_a6_w[1]), 
        .ZN(n2039) );
  OAI221_X1 U1245 ( .B1(n319), .B2(n1693), .C1(n287), .C2(n1694), .A(n2045), 
        .ZN(n2043) );
  AOI22_X1 U1246 ( .A1(n1696), .A2(x7_t2_w[1]), .B1(n1697), .B2(x6_t1_w[1]), 
        .ZN(n2045) );
  OAI221_X1 U1247 ( .B1(n766), .B2(n1668), .C1(n734), .C2(n1669), .A(n1852), 
        .ZN(n1851) );
  AOI22_X1 U1248 ( .A1(n1671), .A2(x17_a7_w[2]), .B1(n1672), .B2(x16_a6_w[2]), 
        .ZN(n1852) );
  OAI221_X1 U1249 ( .B1(n318), .B2(n1693), .C1(n286), .C2(n1694), .A(n1858), 
        .ZN(n1856) );
  AOI22_X1 U1250 ( .A1(n1696), .A2(x7_t2_w[2]), .B1(n1697), .B2(x6_t1_w[2]), 
        .ZN(n1858) );
  OAI221_X1 U1251 ( .B1(n765), .B2(n1668), .C1(n733), .C2(n1669), .A(n1801), 
        .ZN(n1800) );
  AOI22_X1 U1252 ( .A1(n1671), .A2(x17_a7_w[3]), .B1(n1672), .B2(x16_a6_w[3]), 
        .ZN(n1801) );
  OAI221_X1 U1253 ( .B1(n317), .B2(n1693), .C1(n285), .C2(n1694), .A(n1807), 
        .ZN(n1805) );
  AOI22_X1 U1254 ( .A1(n1696), .A2(x7_t2_w[3]), .B1(n1697), .B2(x6_t1_w[3]), 
        .ZN(n1807) );
  OAI221_X1 U1255 ( .B1(n764), .B2(n1668), .C1(n732), .C2(n1669), .A(n1784), 
        .ZN(n1783) );
  AOI22_X1 U1256 ( .A1(n1671), .A2(x17_a7_w[4]), .B1(n1672), .B2(x16_a6_w[4]), 
        .ZN(n1784) );
  OAI221_X1 U1257 ( .B1(n316), .B2(n1693), .C1(n284), .C2(n1694), .A(n1790), 
        .ZN(n1788) );
  AOI22_X1 U1258 ( .A1(n1696), .A2(x7_t2_w[4]), .B1(n1697), .B2(x6_t1_w[4]), 
        .ZN(n1790) );
  OAI221_X1 U1259 ( .B1(n763), .B2(n1668), .C1(n731), .C2(n1669), .A(n1767), 
        .ZN(n1766) );
  AOI22_X1 U1260 ( .A1(n1671), .A2(x17_a7_w[5]), .B1(n1672), .B2(x16_a6_w[5]), 
        .ZN(n1767) );
  OAI221_X1 U1261 ( .B1(n315), .B2(n1693), .C1(n283), .C2(n1694), .A(n1773), 
        .ZN(n1771) );
  AOI22_X1 U1262 ( .A1(n1696), .A2(x7_t2_w[5]), .B1(n1697), .B2(x6_t1_w[5]), 
        .ZN(n1773) );
  OAI221_X1 U1263 ( .B1(n762), .B2(n1668), .C1(n730), .C2(n1669), .A(n1750), 
        .ZN(n1749) );
  AOI22_X1 U1264 ( .A1(n1671), .A2(x17_a7_w[6]), .B1(n1672), .B2(x16_a6_w[6]), 
        .ZN(n1750) );
  OAI221_X1 U1265 ( .B1(n314), .B2(n1693), .C1(n282), .C2(n1694), .A(n1756), 
        .ZN(n1754) );
  AOI22_X1 U1266 ( .A1(n1696), .A2(x7_t2_w[6]), .B1(n1697), .B2(x6_t1_w[6]), 
        .ZN(n1756) );
  OAI221_X1 U1267 ( .B1(n761), .B2(n1668), .C1(n729), .C2(n1669), .A(n1733), 
        .ZN(n1732) );
  AOI22_X1 U1268 ( .A1(n1671), .A2(x17_a7_w[7]), .B1(n1672), .B2(x16_a6_w[7]), 
        .ZN(n1733) );
  OAI221_X1 U1269 ( .B1(n313), .B2(n1693), .C1(n281), .C2(n1694), .A(n1739), 
        .ZN(n1737) );
  AOI22_X1 U1270 ( .A1(n1696), .A2(x7_t2_w[7]), .B1(n1697), .B2(x6_t1_w[7]), 
        .ZN(n1739) );
  OAI221_X1 U1271 ( .B1(n760), .B2(n1668), .C1(n728), .C2(n1669), .A(n1716), 
        .ZN(n1715) );
  AOI22_X1 U1272 ( .A1(n1671), .A2(x17_a7_w[8]), .B1(n1672), .B2(x16_a6_w[8]), 
        .ZN(n1716) );
  OAI221_X1 U1273 ( .B1(n312), .B2(n1693), .C1(n280), .C2(n1694), .A(n1722), 
        .ZN(n1720) );
  AOI22_X1 U1274 ( .A1(n1696), .A2(x7_t2_w[8]), .B1(n1697), .B2(x6_t1_w[8]), 
        .ZN(n1722) );
  OAI221_X1 U1275 ( .B1(n759), .B2(n1668), .C1(n727), .C2(n1669), .A(n1670), 
        .ZN(n1667) );
  AOI22_X1 U1276 ( .A1(n1671), .A2(x17_a7_w[9]), .B1(n1672), .B2(x16_a6_w[9]), 
        .ZN(n1670) );
  OAI221_X1 U1277 ( .B1(n311), .B2(n1693), .C1(n279), .C2(n1694), .A(n1695), 
        .ZN(n1689) );
  AOI22_X1 U1278 ( .A1(n1696), .A2(x7_t2_w[9]), .B1(n1697), .B2(x6_t1_w[9]), 
        .ZN(n1695) );
  OAI221_X1 U1279 ( .B1(n758), .B2(n1668), .C1(n726), .C2(n1669), .A(n2209), 
        .ZN(n2208) );
  AOI22_X1 U1280 ( .A1(n1671), .A2(x17_a7_w[10]), .B1(n1672), .B2(x16_a6_w[10]), .ZN(n2209) );
  OAI221_X1 U1281 ( .B1(n310), .B2(n1693), .C1(n278), .C2(n1694), .A(n2215), 
        .ZN(n2213) );
  AOI22_X1 U1282 ( .A1(n1696), .A2(x7_t2_w[10]), .B1(n1697), .B2(x6_t1_w[10]), 
        .ZN(n2215) );
  OAI221_X1 U1283 ( .B1(n757), .B2(n1668), .C1(n725), .C2(n1669), .A(n2192), 
        .ZN(n2191) );
  AOI22_X1 U1284 ( .A1(n1671), .A2(x17_a7_w[11]), .B1(n1672), .B2(x16_a6_w[11]), .ZN(n2192) );
  OAI221_X1 U1285 ( .B1(n309), .B2(n1693), .C1(n277), .C2(n1694), .A(n2198), 
        .ZN(n2196) );
  AOI22_X1 U1286 ( .A1(n1696), .A2(x7_t2_w[11]), .B1(n1697), .B2(x6_t1_w[11]), 
        .ZN(n2198) );
  OAI221_X1 U1287 ( .B1(n756), .B2(n1668), .C1(n724), .C2(n1669), .A(n2175), 
        .ZN(n2174) );
  AOI22_X1 U1288 ( .A1(n1671), .A2(x17_a7_w[12]), .B1(n1672), .B2(x16_a6_w[12]), .ZN(n2175) );
  OAI221_X1 U1289 ( .B1(n308), .B2(n1693), .C1(n276), .C2(n1694), .A(n2181), 
        .ZN(n2179) );
  AOI22_X1 U1290 ( .A1(n1696), .A2(x7_t2_w[12]), .B1(n1697), .B2(x6_t1_w[12]), 
        .ZN(n2181) );
  OAI221_X1 U1291 ( .B1(n755), .B2(n1668), .C1(n723), .C2(n1669), .A(n2158), 
        .ZN(n2157) );
  AOI22_X1 U1292 ( .A1(n1671), .A2(x17_a7_w[13]), .B1(n1672), .B2(x16_a6_w[13]), .ZN(n2158) );
  OAI221_X1 U1293 ( .B1(n307), .B2(n1693), .C1(n275), .C2(n1694), .A(n2164), 
        .ZN(n2162) );
  AOI22_X1 U1294 ( .A1(n1696), .A2(x7_t2_w[13]), .B1(n1697), .B2(x6_t1_w[13]), 
        .ZN(n2164) );
  OAI221_X1 U1295 ( .B1(n754), .B2(n1668), .C1(n722), .C2(n1669), .A(n2141), 
        .ZN(n2140) );
  AOI22_X1 U1296 ( .A1(n1671), .A2(x17_a7_w[14]), .B1(n1672), .B2(x16_a6_w[14]), .ZN(n2141) );
  OAI221_X1 U1297 ( .B1(n306), .B2(n1693), .C1(n274), .C2(n1694), .A(n2147), 
        .ZN(n2145) );
  AOI22_X1 U1298 ( .A1(n1696), .A2(x7_t2_w[14]), .B1(n1697), .B2(x6_t1_w[14]), 
        .ZN(n2147) );
  OAI221_X1 U1299 ( .B1(n753), .B2(n1668), .C1(n721), .C2(n1669), .A(n2124), 
        .ZN(n2123) );
  AOI22_X1 U1300 ( .A1(n1671), .A2(x17_a7_w[15]), .B1(n1672), .B2(x16_a6_w[15]), .ZN(n2124) );
  OAI221_X1 U1301 ( .B1(n305), .B2(n1693), .C1(n273), .C2(n1694), .A(n2130), 
        .ZN(n2128) );
  AOI22_X1 U1302 ( .A1(n1696), .A2(x7_t2_w[15]), .B1(n1697), .B2(x6_t1_w[15]), 
        .ZN(n2130) );
  OAI221_X1 U1303 ( .B1(n752), .B2(n1668), .C1(n720), .C2(n1669), .A(n2107), 
        .ZN(n2106) );
  AOI22_X1 U1304 ( .A1(n1671), .A2(x17_a7_w[16]), .B1(n1672), .B2(x16_a6_w[16]), .ZN(n2107) );
  OAI221_X1 U1305 ( .B1(n304), .B2(n1693), .C1(n272), .C2(n1694), .A(n2113), 
        .ZN(n2111) );
  AOI22_X1 U1306 ( .A1(n1696), .A2(x7_t2_w[16]), .B1(n1697), .B2(x6_t1_w[16]), 
        .ZN(n2113) );
  OAI221_X1 U1307 ( .B1(n751), .B2(n1668), .C1(n719), .C2(n1669), .A(n2090), 
        .ZN(n2089) );
  AOI22_X1 U1308 ( .A1(n1671), .A2(x17_a7_w[17]), .B1(n1672), .B2(x16_a6_w[17]), .ZN(n2090) );
  OAI221_X1 U1309 ( .B1(n303), .B2(n1693), .C1(n271), .C2(n1694), .A(n2096), 
        .ZN(n2094) );
  AOI22_X1 U1310 ( .A1(n1696), .A2(x7_t2_w[17]), .B1(n1697), .B2(x6_t1_w[17]), 
        .ZN(n2096) );
  OAI221_X1 U1311 ( .B1(n750), .B2(n1668), .C1(n718), .C2(n1669), .A(n2073), 
        .ZN(n2072) );
  AOI22_X1 U1312 ( .A1(n1671), .A2(x17_a7_w[18]), .B1(n1672), .B2(x16_a6_w[18]), .ZN(n2073) );
  OAI221_X1 U1313 ( .B1(n302), .B2(n1693), .C1(n270), .C2(n1694), .A(n2079), 
        .ZN(n2077) );
  AOI22_X1 U1314 ( .A1(n1696), .A2(x7_t2_w[18]), .B1(n1697), .B2(x6_t1_w[18]), 
        .ZN(n2079) );
  OAI221_X1 U1315 ( .B1(n749), .B2(n1668), .C1(n717), .C2(n1669), .A(n2056), 
        .ZN(n2055) );
  AOI22_X1 U1316 ( .A1(n1671), .A2(x17_a7_w[19]), .B1(n1672), .B2(x16_a6_w[19]), .ZN(n2056) );
  OAI221_X1 U1317 ( .B1(n301), .B2(n1693), .C1(n269), .C2(n1694), .A(n2062), 
        .ZN(n2060) );
  AOI22_X1 U1318 ( .A1(n1696), .A2(x7_t2_w[19]), .B1(n1697), .B2(x6_t1_w[19]), 
        .ZN(n2062) );
  OAI221_X1 U1319 ( .B1(n748), .B2(n1668), .C1(n716), .C2(n1669), .A(n2022), 
        .ZN(n2021) );
  AOI22_X1 U1320 ( .A1(n1671), .A2(x17_a7_w[20]), .B1(n1672), .B2(x16_a6_w[20]), .ZN(n2022) );
  OAI221_X1 U1321 ( .B1(n300), .B2(n1693), .C1(n268), .C2(n1694), .A(n2028), 
        .ZN(n2026) );
  AOI22_X1 U1322 ( .A1(n1696), .A2(x7_t2_w[20]), .B1(n1697), .B2(x6_t1_w[20]), 
        .ZN(n2028) );
  OAI221_X1 U1323 ( .B1(n747), .B2(n1668), .C1(n715), .C2(n1669), .A(n2005), 
        .ZN(n2004) );
  AOI22_X1 U1324 ( .A1(n1671), .A2(x17_a7_w[21]), .B1(n1672), .B2(x16_a6_w[21]), .ZN(n2005) );
  OAI221_X1 U1325 ( .B1(n299), .B2(n1693), .C1(n267), .C2(n1694), .A(n2011), 
        .ZN(n2009) );
  AOI22_X1 U1326 ( .A1(n1696), .A2(x7_t2_w[21]), .B1(n1697), .B2(x6_t1_w[21]), 
        .ZN(n2011) );
  OAI221_X1 U1327 ( .B1(n746), .B2(n1668), .C1(n714), .C2(n1669), .A(n1988), 
        .ZN(n1987) );
  AOI22_X1 U1328 ( .A1(n1671), .A2(x17_a7_w[22]), .B1(n1672), .B2(x16_a6_w[22]), .ZN(n1988) );
  OAI221_X1 U1329 ( .B1(n298), .B2(n1693), .C1(n266), .C2(n1694), .A(n1994), 
        .ZN(n1992) );
  AOI22_X1 U1330 ( .A1(n1696), .A2(x7_t2_w[22]), .B1(n1697), .B2(x6_t1_w[22]), 
        .ZN(n1994) );
  OAI221_X1 U1331 ( .B1(n745), .B2(n1668), .C1(n713), .C2(n1669), .A(n1971), 
        .ZN(n1970) );
  AOI22_X1 U1332 ( .A1(n1671), .A2(x17_a7_w[23]), .B1(n1672), .B2(x16_a6_w[23]), .ZN(n1971) );
  OAI221_X1 U1333 ( .B1(n297), .B2(n1693), .C1(n265), .C2(n1694), .A(n1977), 
        .ZN(n1975) );
  AOI22_X1 U1334 ( .A1(n1696), .A2(x7_t2_w[23]), .B1(n1697), .B2(x6_t1_w[23]), 
        .ZN(n1977) );
  OAI221_X1 U1335 ( .B1(n744), .B2(n1668), .C1(n712), .C2(n1669), .A(n1954), 
        .ZN(n1953) );
  AOI22_X1 U1336 ( .A1(n1671), .A2(x17_a7_w[24]), .B1(n1672), .B2(x16_a6_w[24]), .ZN(n1954) );
  OAI221_X1 U1337 ( .B1(n296), .B2(n1693), .C1(n264), .C2(n1694), .A(n1960), 
        .ZN(n1958) );
  AOI22_X1 U1338 ( .A1(n1696), .A2(x7_t2_w[24]), .B1(n1697), .B2(x6_t1_w[24]), 
        .ZN(n1960) );
  OAI221_X1 U1339 ( .B1(n743), .B2(n1668), .C1(n711), .C2(n1669), .A(n1937), 
        .ZN(n1936) );
  AOI22_X1 U1340 ( .A1(n1671), .A2(x17_a7_w[25]), .B1(n1672), .B2(x16_a6_w[25]), .ZN(n1937) );
  OAI221_X1 U1341 ( .B1(n295), .B2(n1693), .C1(n263), .C2(n1694), .A(n1943), 
        .ZN(n1941) );
  AOI22_X1 U1342 ( .A1(n1696), .A2(x7_t2_w[25]), .B1(n1697), .B2(x6_t1_w[25]), 
        .ZN(n1943) );
  OAI221_X1 U1343 ( .B1(n742), .B2(n1668), .C1(n710), .C2(n1669), .A(n1920), 
        .ZN(n1919) );
  AOI22_X1 U1344 ( .A1(n1671), .A2(x17_a7_w[26]), .B1(n1672), .B2(x16_a6_w[26]), .ZN(n1920) );
  OAI221_X1 U1345 ( .B1(n294), .B2(n1693), .C1(n262), .C2(n1694), .A(n1926), 
        .ZN(n1924) );
  AOI22_X1 U1346 ( .A1(n1696), .A2(x7_t2_w[26]), .B1(n1697), .B2(x6_t1_w[26]), 
        .ZN(n1926) );
  OAI221_X1 U1347 ( .B1(n741), .B2(n1668), .C1(n709), .C2(n1669), .A(n1903), 
        .ZN(n1902) );
  AOI22_X1 U1348 ( .A1(n1671), .A2(x17_a7_w[27]), .B1(n1672), .B2(x16_a6_w[27]), .ZN(n1903) );
  OAI221_X1 U1349 ( .B1(n293), .B2(n1693), .C1(n261), .C2(n1694), .A(n1909), 
        .ZN(n1907) );
  AOI22_X1 U1350 ( .A1(n1696), .A2(x7_t2_w[27]), .B1(n1697), .B2(x6_t1_w[27]), 
        .ZN(n1909) );
  OAI221_X1 U1351 ( .B1(n740), .B2(n1668), .C1(n708), .C2(n1669), .A(n1886), 
        .ZN(n1885) );
  AOI22_X1 U1352 ( .A1(n1671), .A2(x17_a7_w[28]), .B1(n1672), .B2(x16_a6_w[28]), .ZN(n1886) );
  OAI221_X1 U1353 ( .B1(n292), .B2(n1693), .C1(n260), .C2(n1694), .A(n1892), 
        .ZN(n1890) );
  AOI22_X1 U1354 ( .A1(n1696), .A2(x7_t2_w[28]), .B1(n1697), .B2(x6_t1_w[28]), 
        .ZN(n1892) );
  OAI221_X1 U1355 ( .B1(n739), .B2(n1668), .C1(n707), .C2(n1669), .A(n1869), 
        .ZN(n1868) );
  AOI22_X1 U1356 ( .A1(n1671), .A2(x17_a7_w[29]), .B1(n1672), .B2(x16_a6_w[29]), .ZN(n1869) );
  OAI221_X1 U1357 ( .B1(n291), .B2(n1693), .C1(n259), .C2(n1694), .A(n1875), 
        .ZN(n1873) );
  AOI22_X1 U1358 ( .A1(n1696), .A2(x7_t2_w[29]), .B1(n1697), .B2(x6_t1_w[29]), 
        .ZN(n1875) );
  OAI221_X1 U1359 ( .B1(n738), .B2(n1668), .C1(n706), .C2(n1669), .A(n1835), 
        .ZN(n1834) );
  AOI22_X1 U1360 ( .A1(n1671), .A2(x17_a7_w[30]), .B1(n1672), .B2(x16_a6_w[30]), .ZN(n1835) );
  OAI221_X1 U1361 ( .B1(n290), .B2(n1693), .C1(n258), .C2(n1694), .A(n1841), 
        .ZN(n1839) );
  AOI22_X1 U1362 ( .A1(n1696), .A2(x7_t2_w[30]), .B1(n1697), .B2(x6_t1_w[30]), 
        .ZN(n1841) );
  OAI221_X1 U1363 ( .B1(n737), .B2(n1668), .C1(n705), .C2(n1669), .A(n1818), 
        .ZN(n1817) );
  AOI22_X1 U1364 ( .A1(n1671), .A2(x17_a7_w[31]), .B1(n1672), .B2(x16_a6_w[31]), .ZN(n1818) );
  OAI221_X1 U1365 ( .B1(n289), .B2(n1693), .C1(n257), .C2(n1694), .A(n1824), 
        .ZN(n1822) );
  AOI22_X1 U1366 ( .A1(n1696), .A2(x7_t2_w[31]), .B1(n1697), .B2(x6_t1_w[31]), 
        .ZN(n1824) );
  OAI22_X1 U1367 ( .A1(n3695), .A2(n599), .B1(n70), .B2(n960), .ZN(n2779) );
  OAI22_X1 U1368 ( .A1(n3679), .A2(n598), .B1(n70), .B2(n959), .ZN(n2780) );
  OAI22_X1 U1369 ( .A1(n3663), .A2(n599), .B1(n70), .B2(n958), .ZN(n2781) );
  OAI22_X1 U1370 ( .A1(n3647), .A2(n598), .B1(n70), .B2(n957), .ZN(n2782) );
  OAI22_X1 U1371 ( .A1(n3631), .A2(n599), .B1(n70), .B2(n956), .ZN(n2783) );
  OAI22_X1 U1372 ( .A1(n3615), .A2(n598), .B1(n70), .B2(n955), .ZN(n2784) );
  OAI22_X1 U1373 ( .A1(n3599), .A2(n599), .B1(n70), .B2(n954), .ZN(n2785) );
  OAI22_X1 U1374 ( .A1(n3583), .A2(n598), .B1(n70), .B2(n953), .ZN(n2786) );
  OAI22_X1 U1375 ( .A1(n3567), .A2(n599), .B1(n70), .B2(n952), .ZN(n2787) );
  OAI22_X1 U1376 ( .A1(n3551), .A2(n599), .B1(n70), .B2(n951), .ZN(n2788) );
  OAI22_X1 U1377 ( .A1(n3535), .A2(n599), .B1(n70), .B2(n950), .ZN(n2789) );
  OAI22_X1 U1378 ( .A1(n3519), .A2(n599), .B1(n70), .B2(n949), .ZN(n2790) );
  OAI22_X1 U1379 ( .A1(n3503), .A2(n599), .B1(n70), .B2(n948), .ZN(n2791) );
  OAI22_X1 U1380 ( .A1(n3487), .A2(n599), .B1(n70), .B2(n947), .ZN(n2792) );
  OAI22_X1 U1381 ( .A1(n3471), .A2(n599), .B1(n70), .B2(n946), .ZN(n2793) );
  OAI22_X1 U1382 ( .A1(n3455), .A2(n599), .B1(n70), .B2(n945), .ZN(n2794) );
  OAI22_X1 U1383 ( .A1(n3439), .A2(n599), .B1(n70), .B2(n944), .ZN(n2795) );
  OAI22_X1 U1384 ( .A1(n3423), .A2(n599), .B1(n70), .B2(n943), .ZN(n2796) );
  OAI22_X1 U1385 ( .A1(n3407), .A2(n599), .B1(n70), .B2(n942), .ZN(n2797) );
  OAI22_X1 U1386 ( .A1(n3391), .A2(n599), .B1(n70), .B2(n941), .ZN(n2798) );
  OAI22_X1 U1387 ( .A1(n3375), .A2(n598), .B1(n70), .B2(n940), .ZN(n2799) );
  OAI22_X1 U1388 ( .A1(n3359), .A2(n598), .B1(n70), .B2(n939), .ZN(n2800) );
  OAI22_X1 U1389 ( .A1(n3343), .A2(n598), .B1(n70), .B2(n938), .ZN(n2801) );
  OAI22_X1 U1390 ( .A1(n3327), .A2(n598), .B1(n70), .B2(n937), .ZN(n2802) );
  OAI22_X1 U1391 ( .A1(n3311), .A2(n598), .B1(n70), .B2(n936), .ZN(n2803) );
  OAI22_X1 U1392 ( .A1(n3295), .A2(n598), .B1(n70), .B2(n935), .ZN(n2804) );
  OAI22_X1 U1393 ( .A1(n2361), .A2(n598), .B1(n70), .B2(n934), .ZN(n2805) );
  OAI22_X1 U1394 ( .A1(n1058), .A2(n598), .B1(n70), .B2(n933), .ZN(n2806) );
  OAI22_X1 U1395 ( .A1(n1042), .A2(n598), .B1(n70), .B2(n932), .ZN(n2807) );
  OAI22_X1 U1396 ( .A1(n1026), .A2(n598), .B1(n70), .B2(n931), .ZN(n2808) );
  OAI22_X1 U1397 ( .A1(n1010), .A2(n598), .B1(n70), .B2(n930), .ZN(n2809) );
  OAI22_X1 U1398 ( .A1(n994), .A2(n598), .B1(n70), .B2(n929), .ZN(n2810) );
  OAI22_X1 U1399 ( .A1(n3695), .A2(n590), .B1(n69), .B2(n928), .ZN(n2811) );
  OAI22_X1 U1400 ( .A1(n3679), .A2(n589), .B1(n69), .B2(n927), .ZN(n2812) );
  OAI22_X1 U1401 ( .A1(n3663), .A2(n590), .B1(n69), .B2(n926), .ZN(n2813) );
  OAI22_X1 U1402 ( .A1(n3647), .A2(n589), .B1(n69), .B2(n925), .ZN(n2814) );
  OAI22_X1 U1403 ( .A1(n3631), .A2(n590), .B1(n69), .B2(n924), .ZN(n2815) );
  OAI22_X1 U1404 ( .A1(n3615), .A2(n589), .B1(n69), .B2(n923), .ZN(n2816) );
  OAI22_X1 U1405 ( .A1(n3599), .A2(n590), .B1(n69), .B2(n922), .ZN(n2817) );
  OAI22_X1 U1406 ( .A1(n3583), .A2(n589), .B1(n69), .B2(n921), .ZN(n2818) );
  OAI22_X1 U1407 ( .A1(n3567), .A2(n590), .B1(n69), .B2(n920), .ZN(n2819) );
  OAI22_X1 U1408 ( .A1(n3551), .A2(n590), .B1(n69), .B2(n919), .ZN(n2820) );
  OAI22_X1 U1409 ( .A1(n3535), .A2(n590), .B1(n69), .B2(n918), .ZN(n2821) );
  OAI22_X1 U1410 ( .A1(n3519), .A2(n590), .B1(n69), .B2(n917), .ZN(n2822) );
  OAI22_X1 U1411 ( .A1(n3503), .A2(n590), .B1(n69), .B2(n916), .ZN(n2823) );
  OAI22_X1 U1412 ( .A1(n3487), .A2(n590), .B1(n69), .B2(n915), .ZN(n2824) );
  OAI22_X1 U1413 ( .A1(n3471), .A2(n590), .B1(n69), .B2(n914), .ZN(n2825) );
  OAI22_X1 U1414 ( .A1(n3455), .A2(n590), .B1(n69), .B2(n913), .ZN(n2826) );
  OAI22_X1 U1415 ( .A1(n3439), .A2(n590), .B1(n69), .B2(n912), .ZN(n2827) );
  OAI22_X1 U1416 ( .A1(n3423), .A2(n590), .B1(n69), .B2(n911), .ZN(n2828) );
  OAI22_X1 U1417 ( .A1(n3407), .A2(n590), .B1(n69), .B2(n910), .ZN(n2829) );
  OAI22_X1 U1418 ( .A1(n3391), .A2(n590), .B1(n69), .B2(n909), .ZN(n2830) );
  OAI22_X1 U1419 ( .A1(n3375), .A2(n589), .B1(n69), .B2(n908), .ZN(n2831) );
  OAI22_X1 U1420 ( .A1(n3359), .A2(n589), .B1(n69), .B2(n907), .ZN(n2832) );
  OAI22_X1 U1421 ( .A1(n3343), .A2(n589), .B1(n69), .B2(n906), .ZN(n2833) );
  OAI22_X1 U1422 ( .A1(n3327), .A2(n589), .B1(n69), .B2(n905), .ZN(n2834) );
  OAI22_X1 U1423 ( .A1(n3311), .A2(n589), .B1(n69), .B2(n904), .ZN(n2835) );
  OAI22_X1 U1424 ( .A1(n3295), .A2(n589), .B1(n69), .B2(n903), .ZN(n2836) );
  OAI22_X1 U1425 ( .A1(n2361), .A2(n589), .B1(n69), .B2(n902), .ZN(n2837) );
  OAI22_X1 U1426 ( .A1(n1058), .A2(n589), .B1(n69), .B2(n901), .ZN(n2838) );
  OAI22_X1 U1427 ( .A1(n1042), .A2(n589), .B1(n69), .B2(n900), .ZN(n2839) );
  OAI22_X1 U1428 ( .A1(n1026), .A2(n589), .B1(n69), .B2(n899), .ZN(n2840) );
  OAI22_X1 U1429 ( .A1(n1010), .A2(n589), .B1(n69), .B2(n898), .ZN(n2841) );
  OAI22_X1 U1430 ( .A1(n994), .A2(n589), .B1(n69), .B2(n897), .ZN(n2842) );
  OAI22_X1 U1431 ( .A1(n3695), .A2(n435), .B1(n71), .B2(n832), .ZN(n2843) );
  OAI22_X1 U1432 ( .A1(n3679), .A2(n434), .B1(n71), .B2(n831), .ZN(n2844) );
  OAI22_X1 U1433 ( .A1(n3663), .A2(n435), .B1(n71), .B2(n830), .ZN(n2845) );
  OAI22_X1 U1434 ( .A1(n3647), .A2(n434), .B1(n71), .B2(n829), .ZN(n2846) );
  OAI22_X1 U1435 ( .A1(n3631), .A2(n435), .B1(n71), .B2(n828), .ZN(n2847) );
  OAI22_X1 U1436 ( .A1(n3615), .A2(n434), .B1(n71), .B2(n827), .ZN(n2848) );
  OAI22_X1 U1437 ( .A1(n3599), .A2(n435), .B1(n71), .B2(n826), .ZN(n2849) );
  OAI22_X1 U1438 ( .A1(n3583), .A2(n434), .B1(n71), .B2(n825), .ZN(n2850) );
  OAI22_X1 U1439 ( .A1(n3567), .A2(n435), .B1(n71), .B2(n824), .ZN(n2851) );
  OAI22_X1 U1440 ( .A1(n3551), .A2(n435), .B1(n71), .B2(n823), .ZN(n2852) );
  OAI22_X1 U1441 ( .A1(n3535), .A2(n435), .B1(n71), .B2(n822), .ZN(n2853) );
  OAI22_X1 U1442 ( .A1(n3519), .A2(n435), .B1(n71), .B2(n821), .ZN(n2854) );
  OAI22_X1 U1443 ( .A1(n3503), .A2(n435), .B1(n71), .B2(n820), .ZN(n2855) );
  OAI22_X1 U1444 ( .A1(n3487), .A2(n435), .B1(n71), .B2(n819), .ZN(n2856) );
  OAI22_X1 U1445 ( .A1(n3471), .A2(n435), .B1(n71), .B2(n818), .ZN(n2857) );
  OAI22_X1 U1446 ( .A1(n3455), .A2(n435), .B1(n71), .B2(n817), .ZN(n2858) );
  OAI22_X1 U1447 ( .A1(n3439), .A2(n435), .B1(n71), .B2(n816), .ZN(n2859) );
  OAI22_X1 U1448 ( .A1(n3423), .A2(n435), .B1(n71), .B2(n815), .ZN(n2860) );
  OAI22_X1 U1449 ( .A1(n3407), .A2(n435), .B1(n71), .B2(n814), .ZN(n2861) );
  OAI22_X1 U1450 ( .A1(n3391), .A2(n435), .B1(n71), .B2(n813), .ZN(n2862) );
  OAI22_X1 U1451 ( .A1(n3375), .A2(n434), .B1(n71), .B2(n812), .ZN(n2863) );
  OAI22_X1 U1452 ( .A1(n3359), .A2(n434), .B1(n71), .B2(n811), .ZN(n2864) );
  OAI22_X1 U1453 ( .A1(n3343), .A2(n434), .B1(n71), .B2(n810), .ZN(n2865) );
  OAI22_X1 U1454 ( .A1(n3327), .A2(n434), .B1(n71), .B2(n809), .ZN(n2866) );
  OAI22_X1 U1455 ( .A1(n3311), .A2(n434), .B1(n71), .B2(n808), .ZN(n2867) );
  OAI22_X1 U1456 ( .A1(n3295), .A2(n434), .B1(n71), .B2(n807), .ZN(n2868) );
  OAI22_X1 U1457 ( .A1(n2361), .A2(n434), .B1(n71), .B2(n806), .ZN(n2869) );
  OAI22_X1 U1458 ( .A1(n1058), .A2(n434), .B1(n71), .B2(n805), .ZN(n2870) );
  OAI22_X1 U1459 ( .A1(n1042), .A2(n434), .B1(n71), .B2(n804), .ZN(n2871) );
  OAI22_X1 U1460 ( .A1(n1026), .A2(n434), .B1(n71), .B2(n803), .ZN(n2872) );
  OAI22_X1 U1461 ( .A1(n1010), .A2(n434), .B1(n71), .B2(n802), .ZN(n2873) );
  OAI22_X1 U1462 ( .A1(n994), .A2(n434), .B1(n71), .B2(n801), .ZN(n2874) );
  OAI22_X1 U1463 ( .A1(n3695), .A2(n426), .B1(n78), .B2(n800), .ZN(n2875) );
  OAI22_X1 U1464 ( .A1(n3679), .A2(n425), .B1(n78), .B2(n799), .ZN(n2876) );
  OAI22_X1 U1465 ( .A1(n3663), .A2(n426), .B1(n78), .B2(n798), .ZN(n2877) );
  OAI22_X1 U1466 ( .A1(n3647), .A2(n425), .B1(n78), .B2(n797), .ZN(n2878) );
  OAI22_X1 U1467 ( .A1(n3631), .A2(n426), .B1(n78), .B2(n796), .ZN(n2879) );
  OAI22_X1 U1468 ( .A1(n3615), .A2(n425), .B1(n78), .B2(n795), .ZN(n2880) );
  OAI22_X1 U1469 ( .A1(n3599), .A2(n426), .B1(n78), .B2(n794), .ZN(n2881) );
  OAI22_X1 U1470 ( .A1(n3583), .A2(n425), .B1(n78), .B2(n793), .ZN(n2882) );
  OAI22_X1 U1471 ( .A1(n3567), .A2(n426), .B1(n78), .B2(n792), .ZN(n2883) );
  OAI22_X1 U1472 ( .A1(n3551), .A2(n426), .B1(n78), .B2(n791), .ZN(n2884) );
  OAI22_X1 U1473 ( .A1(n3535), .A2(n426), .B1(n78), .B2(n790), .ZN(n2885) );
  OAI22_X1 U1474 ( .A1(n3519), .A2(n426), .B1(n78), .B2(n789), .ZN(n2886) );
  OAI22_X1 U1475 ( .A1(n3503), .A2(n426), .B1(n78), .B2(n788), .ZN(n2887) );
  OAI22_X1 U1476 ( .A1(n3487), .A2(n426), .B1(n78), .B2(n787), .ZN(n2888) );
  OAI22_X1 U1477 ( .A1(n3471), .A2(n426), .B1(n78), .B2(n786), .ZN(n2889) );
  OAI22_X1 U1478 ( .A1(n3455), .A2(n426), .B1(n78), .B2(n785), .ZN(n2890) );
  OAI22_X1 U1479 ( .A1(n3439), .A2(n426), .B1(n78), .B2(n784), .ZN(n2891) );
  OAI22_X1 U1480 ( .A1(n3423), .A2(n426), .B1(n78), .B2(n783), .ZN(n2892) );
  OAI22_X1 U1481 ( .A1(n3407), .A2(n426), .B1(n78), .B2(n782), .ZN(n2893) );
  OAI22_X1 U1482 ( .A1(n3391), .A2(n426), .B1(n78), .B2(n781), .ZN(n2894) );
  OAI22_X1 U1483 ( .A1(n3375), .A2(n425), .B1(n78), .B2(n780), .ZN(n2895) );
  OAI22_X1 U1484 ( .A1(n3359), .A2(n425), .B1(n78), .B2(n779), .ZN(n2896) );
  OAI22_X1 U1485 ( .A1(n3343), .A2(n425), .B1(n78), .B2(n778), .ZN(n2897) );
  OAI22_X1 U1486 ( .A1(n3327), .A2(n425), .B1(n78), .B2(n777), .ZN(n2898) );
  OAI22_X1 U1487 ( .A1(n3311), .A2(n425), .B1(n78), .B2(n776), .ZN(n2899) );
  OAI22_X1 U1488 ( .A1(n3295), .A2(n425), .B1(n78), .B2(n775), .ZN(n2900) );
  OAI22_X1 U1489 ( .A1(n2361), .A2(n425), .B1(n78), .B2(n774), .ZN(n2901) );
  OAI22_X1 U1490 ( .A1(n1058), .A2(n425), .B1(n78), .B2(n773), .ZN(n2902) );
  OAI22_X1 U1491 ( .A1(n1042), .A2(n425), .B1(n78), .B2(n772), .ZN(n2903) );
  OAI22_X1 U1492 ( .A1(n1026), .A2(n425), .B1(n78), .B2(n771), .ZN(n2904) );
  OAI22_X1 U1493 ( .A1(n1010), .A2(n425), .B1(n78), .B2(n770), .ZN(n2905) );
  OAI22_X1 U1494 ( .A1(n994), .A2(n425), .B1(n78), .B2(n769), .ZN(n2906) );
  OAI22_X1 U1495 ( .A1(n3695), .A2(n417), .B1(n65), .B2(n768), .ZN(n2907) );
  OAI22_X1 U1496 ( .A1(n3679), .A2(n416), .B1(n65), .B2(n767), .ZN(n2908) );
  OAI22_X1 U1497 ( .A1(n3663), .A2(n417), .B1(n65), .B2(n766), .ZN(n2909) );
  OAI22_X1 U1498 ( .A1(n3647), .A2(n416), .B1(n65), .B2(n765), .ZN(n2910) );
  OAI22_X1 U1499 ( .A1(n3631), .A2(n417), .B1(n65), .B2(n764), .ZN(n2911) );
  OAI22_X1 U1500 ( .A1(n3615), .A2(n416), .B1(n65), .B2(n763), .ZN(n2912) );
  OAI22_X1 U1501 ( .A1(n3599), .A2(n417), .B1(n65), .B2(n762), .ZN(n2913) );
  OAI22_X1 U1502 ( .A1(n3583), .A2(n416), .B1(n65), .B2(n761), .ZN(n2914) );
  OAI22_X1 U1503 ( .A1(n3567), .A2(n417), .B1(n65), .B2(n760), .ZN(n2915) );
  OAI22_X1 U1504 ( .A1(n3551), .A2(n417), .B1(n65), .B2(n759), .ZN(n2916) );
  OAI22_X1 U1505 ( .A1(n3535), .A2(n417), .B1(n65), .B2(n758), .ZN(n2917) );
  OAI22_X1 U1506 ( .A1(n3519), .A2(n417), .B1(n65), .B2(n757), .ZN(n2918) );
  OAI22_X1 U1507 ( .A1(n3503), .A2(n417), .B1(n65), .B2(n756), .ZN(n2919) );
  OAI22_X1 U1508 ( .A1(n3487), .A2(n417), .B1(n65), .B2(n755), .ZN(n2920) );
  OAI22_X1 U1509 ( .A1(n3471), .A2(n417), .B1(n65), .B2(n754), .ZN(n2921) );
  OAI22_X1 U1510 ( .A1(n3455), .A2(n417), .B1(n65), .B2(n753), .ZN(n2922) );
  OAI22_X1 U1511 ( .A1(n3439), .A2(n417), .B1(n65), .B2(n752), .ZN(n2923) );
  OAI22_X1 U1512 ( .A1(n3423), .A2(n417), .B1(n65), .B2(n751), .ZN(n2924) );
  OAI22_X1 U1513 ( .A1(n3407), .A2(n417), .B1(n65), .B2(n750), .ZN(n2925) );
  OAI22_X1 U1514 ( .A1(n3391), .A2(n417), .B1(n65), .B2(n749), .ZN(n2926) );
  OAI22_X1 U1515 ( .A1(n3375), .A2(n416), .B1(n65), .B2(n748), .ZN(n2927) );
  OAI22_X1 U1516 ( .A1(n3359), .A2(n416), .B1(n65), .B2(n747), .ZN(n2928) );
  OAI22_X1 U1517 ( .A1(n3343), .A2(n416), .B1(n65), .B2(n746), .ZN(n2929) );
  OAI22_X1 U1518 ( .A1(n3327), .A2(n416), .B1(n65), .B2(n745), .ZN(n2930) );
  OAI22_X1 U1519 ( .A1(n3311), .A2(n416), .B1(n65), .B2(n744), .ZN(n2931) );
  OAI22_X1 U1520 ( .A1(n3295), .A2(n416), .B1(n65), .B2(n743), .ZN(n2932) );
  OAI22_X1 U1521 ( .A1(n2361), .A2(n416), .B1(n65), .B2(n742), .ZN(n2933) );
  OAI22_X1 U1522 ( .A1(n1058), .A2(n416), .B1(n65), .B2(n741), .ZN(n2934) );
  OAI22_X1 U1523 ( .A1(n1042), .A2(n416), .B1(n65), .B2(n740), .ZN(n2935) );
  OAI22_X1 U1524 ( .A1(n1026), .A2(n416), .B1(n65), .B2(n739), .ZN(n2936) );
  OAI22_X1 U1525 ( .A1(n1010), .A2(n416), .B1(n65), .B2(n738), .ZN(n2937) );
  OAI22_X1 U1526 ( .A1(n994), .A2(n416), .B1(n65), .B2(n737), .ZN(n2938) );
  OAI22_X1 U1527 ( .A1(n3695), .A2(n408), .B1(n72), .B2(n736), .ZN(n2939) );
  OAI22_X1 U1528 ( .A1(n3679), .A2(n407), .B1(n72), .B2(n735), .ZN(n2940) );
  OAI22_X1 U1529 ( .A1(n3663), .A2(n408), .B1(n72), .B2(n734), .ZN(n2941) );
  OAI22_X1 U1530 ( .A1(n3647), .A2(n407), .B1(n72), .B2(n733), .ZN(n2942) );
  OAI22_X1 U1531 ( .A1(n3631), .A2(n408), .B1(n72), .B2(n732), .ZN(n2943) );
  OAI22_X1 U1532 ( .A1(n3615), .A2(n407), .B1(n72), .B2(n731), .ZN(n2944) );
  OAI22_X1 U1533 ( .A1(n3599), .A2(n408), .B1(n72), .B2(n730), .ZN(n2945) );
  OAI22_X1 U1534 ( .A1(n3583), .A2(n407), .B1(n72), .B2(n729), .ZN(n2946) );
  OAI22_X1 U1535 ( .A1(n3567), .A2(n408), .B1(n72), .B2(n728), .ZN(n2947) );
  OAI22_X1 U1536 ( .A1(n3551), .A2(n408), .B1(n72), .B2(n727), .ZN(n2948) );
  OAI22_X1 U1537 ( .A1(n3535), .A2(n408), .B1(n72), .B2(n726), .ZN(n2949) );
  OAI22_X1 U1538 ( .A1(n3519), .A2(n408), .B1(n72), .B2(n725), .ZN(n2950) );
  OAI22_X1 U1539 ( .A1(n3503), .A2(n408), .B1(n72), .B2(n724), .ZN(n2951) );
  OAI22_X1 U1540 ( .A1(n3487), .A2(n408), .B1(n72), .B2(n723), .ZN(n2952) );
  OAI22_X1 U1541 ( .A1(n3471), .A2(n408), .B1(n72), .B2(n722), .ZN(n2953) );
  OAI22_X1 U1542 ( .A1(n3455), .A2(n408), .B1(n72), .B2(n721), .ZN(n2954) );
  OAI22_X1 U1543 ( .A1(n3439), .A2(n408), .B1(n72), .B2(n720), .ZN(n2955) );
  OAI22_X1 U1544 ( .A1(n3423), .A2(n408), .B1(n72), .B2(n719), .ZN(n2956) );
  OAI22_X1 U1545 ( .A1(n3407), .A2(n408), .B1(n72), .B2(n718), .ZN(n2957) );
  OAI22_X1 U1546 ( .A1(n3391), .A2(n408), .B1(n72), .B2(n717), .ZN(n2958) );
  OAI22_X1 U1547 ( .A1(n3375), .A2(n407), .B1(n72), .B2(n716), .ZN(n2959) );
  OAI22_X1 U1548 ( .A1(n3359), .A2(n407), .B1(n72), .B2(n715), .ZN(n2960) );
  OAI22_X1 U1549 ( .A1(n3343), .A2(n407), .B1(n72), .B2(n714), .ZN(n2961) );
  OAI22_X1 U1550 ( .A1(n3327), .A2(n407), .B1(n72), .B2(n713), .ZN(n2962) );
  OAI22_X1 U1551 ( .A1(n3311), .A2(n407), .B1(n72), .B2(n712), .ZN(n2963) );
  OAI22_X1 U1552 ( .A1(n3295), .A2(n407), .B1(n72), .B2(n711), .ZN(n2964) );
  OAI22_X1 U1553 ( .A1(n2361), .A2(n407), .B1(n72), .B2(n710), .ZN(n2965) );
  OAI22_X1 U1554 ( .A1(n1058), .A2(n407), .B1(n72), .B2(n709), .ZN(n2966) );
  OAI22_X1 U1555 ( .A1(n1042), .A2(n407), .B1(n72), .B2(n708), .ZN(n2967) );
  OAI22_X1 U1556 ( .A1(n1026), .A2(n407), .B1(n72), .B2(n707), .ZN(n2968) );
  OAI22_X1 U1557 ( .A1(n1010), .A2(n407), .B1(n72), .B2(n706), .ZN(n2969) );
  OAI22_X1 U1558 ( .A1(n994), .A2(n407), .B1(n72), .B2(n705), .ZN(n2970) );
  OAI22_X1 U1559 ( .A1(n3695), .A2(n363), .B1(n73), .B2(n576), .ZN(n2971) );
  OAI22_X1 U1560 ( .A1(n3679), .A2(n362), .B1(n73), .B2(n575), .ZN(n2972) );
  OAI22_X1 U1561 ( .A1(n3663), .A2(n363), .B1(n73), .B2(n574), .ZN(n2973) );
  OAI22_X1 U1562 ( .A1(n3647), .A2(n362), .B1(n73), .B2(n573), .ZN(n2974) );
  OAI22_X1 U1563 ( .A1(n3631), .A2(n363), .B1(n73), .B2(n572), .ZN(n2975) );
  OAI22_X1 U1564 ( .A1(n3615), .A2(n362), .B1(n73), .B2(n571), .ZN(n2976) );
  OAI22_X1 U1565 ( .A1(n3599), .A2(n363), .B1(n73), .B2(n570), .ZN(n2977) );
  OAI22_X1 U1566 ( .A1(n3583), .A2(n362), .B1(n73), .B2(n569), .ZN(n2978) );
  OAI22_X1 U1567 ( .A1(n3567), .A2(n363), .B1(n73), .B2(n568), .ZN(n2979) );
  OAI22_X1 U1568 ( .A1(n3551), .A2(n363), .B1(n73), .B2(n567), .ZN(n2980) );
  OAI22_X1 U1569 ( .A1(n3535), .A2(n363), .B1(n73), .B2(n566), .ZN(n2981) );
  OAI22_X1 U1570 ( .A1(n3519), .A2(n363), .B1(n73), .B2(n565), .ZN(n2982) );
  OAI22_X1 U1571 ( .A1(n3503), .A2(n363), .B1(n73), .B2(n564), .ZN(n2983) );
  OAI22_X1 U1572 ( .A1(n3487), .A2(n363), .B1(n73), .B2(n563), .ZN(n2984) );
  OAI22_X1 U1573 ( .A1(n3471), .A2(n363), .B1(n73), .B2(n562), .ZN(n2985) );
  OAI22_X1 U1574 ( .A1(n3455), .A2(n363), .B1(n73), .B2(n561), .ZN(n2986) );
  OAI22_X1 U1575 ( .A1(n3439), .A2(n363), .B1(n73), .B2(n560), .ZN(n2987) );
  OAI22_X1 U1576 ( .A1(n3423), .A2(n363), .B1(n73), .B2(n559), .ZN(n2988) );
  OAI22_X1 U1577 ( .A1(n3407), .A2(n363), .B1(n73), .B2(n558), .ZN(n2989) );
  OAI22_X1 U1578 ( .A1(n3391), .A2(n363), .B1(n73), .B2(n557), .ZN(n2990) );
  OAI22_X1 U1579 ( .A1(n3375), .A2(n362), .B1(n73), .B2(n556), .ZN(n2991) );
  OAI22_X1 U1580 ( .A1(n3359), .A2(n362), .B1(n73), .B2(n555), .ZN(n2992) );
  OAI22_X1 U1581 ( .A1(n3343), .A2(n362), .B1(n73), .B2(n554), .ZN(n2993) );
  OAI22_X1 U1582 ( .A1(n3327), .A2(n362), .B1(n73), .B2(n553), .ZN(n2994) );
  OAI22_X1 U1583 ( .A1(n3311), .A2(n362), .B1(n73), .B2(n552), .ZN(n2995) );
  OAI22_X1 U1584 ( .A1(n3295), .A2(n362), .B1(n73), .B2(n551), .ZN(n2996) );
  OAI22_X1 U1585 ( .A1(n2361), .A2(n362), .B1(n73), .B2(n550), .ZN(n2997) );
  OAI22_X1 U1586 ( .A1(n1058), .A2(n362), .B1(n73), .B2(n549), .ZN(n2998) );
  OAI22_X1 U1587 ( .A1(n1042), .A2(n362), .B1(n73), .B2(n548), .ZN(n2999) );
  OAI22_X1 U1588 ( .A1(n1026), .A2(n362), .B1(n73), .B2(n547), .ZN(n3000) );
  OAI22_X1 U1589 ( .A1(n1010), .A2(n362), .B1(n73), .B2(n546), .ZN(n3001) );
  OAI22_X1 U1590 ( .A1(n994), .A2(n362), .B1(n73), .B2(n545), .ZN(n3002) );
  OAI22_X1 U1591 ( .A1(n3695), .A2(n354), .B1(n79), .B2(n544), .ZN(n3003) );
  OAI22_X1 U1592 ( .A1(n3679), .A2(n353), .B1(n79), .B2(n543), .ZN(n3004) );
  OAI22_X1 U1593 ( .A1(n3663), .A2(n354), .B1(n79), .B2(n542), .ZN(n3005) );
  OAI22_X1 U1594 ( .A1(n3647), .A2(n353), .B1(n79), .B2(n541), .ZN(n3006) );
  OAI22_X1 U1595 ( .A1(n3631), .A2(n354), .B1(n79), .B2(n540), .ZN(n3007) );
  OAI22_X1 U1596 ( .A1(n3615), .A2(n353), .B1(n79), .B2(n539), .ZN(n3008) );
  OAI22_X1 U1597 ( .A1(n3599), .A2(n354), .B1(n79), .B2(n538), .ZN(n3009) );
  OAI22_X1 U1598 ( .A1(n3583), .A2(n353), .B1(n79), .B2(n537), .ZN(n3010) );
  OAI22_X1 U1599 ( .A1(n3567), .A2(n354), .B1(n79), .B2(n536), .ZN(n3011) );
  OAI22_X1 U1600 ( .A1(n3551), .A2(n354), .B1(n79), .B2(n535), .ZN(n3012) );
  OAI22_X1 U1601 ( .A1(n3535), .A2(n354), .B1(n79), .B2(n534), .ZN(n3013) );
  OAI22_X1 U1602 ( .A1(n3519), .A2(n354), .B1(n79), .B2(n533), .ZN(n3014) );
  OAI22_X1 U1603 ( .A1(n3503), .A2(n354), .B1(n79), .B2(n532), .ZN(n3015) );
  OAI22_X1 U1604 ( .A1(n3487), .A2(n354), .B1(n79), .B2(n531), .ZN(n3016) );
  OAI22_X1 U1605 ( .A1(n3471), .A2(n354), .B1(n79), .B2(n530), .ZN(n3017) );
  OAI22_X1 U1606 ( .A1(n3455), .A2(n354), .B1(n79), .B2(n529), .ZN(n3018) );
  OAI22_X1 U1607 ( .A1(n3439), .A2(n354), .B1(n79), .B2(n528), .ZN(n3019) );
  OAI22_X1 U1608 ( .A1(n3423), .A2(n354), .B1(n79), .B2(n527), .ZN(n3020) );
  OAI22_X1 U1609 ( .A1(n3407), .A2(n354), .B1(n79), .B2(n526), .ZN(n3021) );
  OAI22_X1 U1610 ( .A1(n3391), .A2(n354), .B1(n79), .B2(n525), .ZN(n3022) );
  OAI22_X1 U1611 ( .A1(n3375), .A2(n353), .B1(n79), .B2(n524), .ZN(n3023) );
  OAI22_X1 U1612 ( .A1(n3359), .A2(n353), .B1(n79), .B2(n523), .ZN(n3024) );
  OAI22_X1 U1613 ( .A1(n3343), .A2(n353), .B1(n79), .B2(n522), .ZN(n3025) );
  OAI22_X1 U1614 ( .A1(n3327), .A2(n353), .B1(n79), .B2(n521), .ZN(n3026) );
  OAI22_X1 U1615 ( .A1(n3311), .A2(n353), .B1(n79), .B2(n520), .ZN(n3027) );
  OAI22_X1 U1616 ( .A1(n3295), .A2(n353), .B1(n79), .B2(n519), .ZN(n3028) );
  OAI22_X1 U1617 ( .A1(n2361), .A2(n353), .B1(n79), .B2(n518), .ZN(n3029) );
  OAI22_X1 U1618 ( .A1(n1058), .A2(n353), .B1(n79), .B2(n517), .ZN(n3030) );
  OAI22_X1 U1619 ( .A1(n1042), .A2(n353), .B1(n79), .B2(n516), .ZN(n3031) );
  OAI22_X1 U1620 ( .A1(n1026), .A2(n353), .B1(n79), .B2(n515), .ZN(n3032) );
  OAI22_X1 U1621 ( .A1(n1010), .A2(n353), .B1(n79), .B2(n514), .ZN(n3033) );
  OAI22_X1 U1622 ( .A1(n994), .A2(n353), .B1(n79), .B2(n513), .ZN(n3034) );
  OAI22_X1 U1623 ( .A1(n3695), .A2(n345), .B1(n66), .B2(n512), .ZN(n3035) );
  OAI22_X1 U1624 ( .A1(n3679), .A2(n344), .B1(n66), .B2(n511), .ZN(n3036) );
  OAI22_X1 U1625 ( .A1(n3663), .A2(n345), .B1(n66), .B2(n510), .ZN(n3037) );
  OAI22_X1 U1626 ( .A1(n3647), .A2(n344), .B1(n66), .B2(n509), .ZN(n3038) );
  OAI22_X1 U1627 ( .A1(n3631), .A2(n345), .B1(n66), .B2(n508), .ZN(n3039) );
  OAI22_X1 U1628 ( .A1(n3615), .A2(n344), .B1(n66), .B2(n507), .ZN(n3040) );
  OAI22_X1 U1629 ( .A1(n3599), .A2(n345), .B1(n66), .B2(n506), .ZN(n3041) );
  OAI22_X1 U1630 ( .A1(n3583), .A2(n344), .B1(n66), .B2(n505), .ZN(n3042) );
  OAI22_X1 U1631 ( .A1(n3567), .A2(n345), .B1(n66), .B2(n504), .ZN(n3043) );
  OAI22_X1 U1632 ( .A1(n3551), .A2(n345), .B1(n66), .B2(n503), .ZN(n3044) );
  OAI22_X1 U1633 ( .A1(n3535), .A2(n345), .B1(n66), .B2(n502), .ZN(n3045) );
  OAI22_X1 U1634 ( .A1(n3519), .A2(n345), .B1(n66), .B2(n501), .ZN(n3046) );
  OAI22_X1 U1635 ( .A1(n3503), .A2(n345), .B1(n66), .B2(n500), .ZN(n3047) );
  OAI22_X1 U1636 ( .A1(n3487), .A2(n345), .B1(n66), .B2(n499), .ZN(n3048) );
  OAI22_X1 U1637 ( .A1(n3471), .A2(n345), .B1(n66), .B2(n498), .ZN(n3049) );
  OAI22_X1 U1638 ( .A1(n3455), .A2(n345), .B1(n66), .B2(n497), .ZN(n3050) );
  OAI22_X1 U1639 ( .A1(n3439), .A2(n345), .B1(n66), .B2(n496), .ZN(n3051) );
  OAI22_X1 U1640 ( .A1(n3423), .A2(n345), .B1(n66), .B2(n495), .ZN(n3052) );
  OAI22_X1 U1641 ( .A1(n3407), .A2(n345), .B1(n66), .B2(n494), .ZN(n3053) );
  OAI22_X1 U1642 ( .A1(n3391), .A2(n345), .B1(n66), .B2(n493), .ZN(n3054) );
  OAI22_X1 U1643 ( .A1(n3375), .A2(n344), .B1(n66), .B2(n492), .ZN(n3055) );
  OAI22_X1 U1644 ( .A1(n3359), .A2(n344), .B1(n66), .B2(n491), .ZN(n3056) );
  OAI22_X1 U1645 ( .A1(n3343), .A2(n344), .B1(n66), .B2(n490), .ZN(n3057) );
  OAI22_X1 U1646 ( .A1(n3327), .A2(n344), .B1(n66), .B2(n489), .ZN(n3058) );
  OAI22_X1 U1647 ( .A1(n3311), .A2(n344), .B1(n66), .B2(n488), .ZN(n3059) );
  OAI22_X1 U1648 ( .A1(n3295), .A2(n344), .B1(n66), .B2(n487), .ZN(n3060) );
  OAI22_X1 U1649 ( .A1(n2361), .A2(n344), .B1(n66), .B2(n486), .ZN(n3061) );
  OAI22_X1 U1650 ( .A1(n1058), .A2(n344), .B1(n66), .B2(n485), .ZN(n3062) );
  OAI22_X1 U1651 ( .A1(n1042), .A2(n344), .B1(n66), .B2(n484), .ZN(n3063) );
  OAI22_X1 U1652 ( .A1(n1026), .A2(n344), .B1(n66), .B2(n483), .ZN(n3064) );
  OAI22_X1 U1653 ( .A1(n1010), .A2(n344), .B1(n66), .B2(n482), .ZN(n3065) );
  OAI22_X1 U1654 ( .A1(n994), .A2(n344), .B1(n66), .B2(n481), .ZN(n3066) );
  OAI22_X1 U1655 ( .A1(n3695), .A2(n336), .B1(n74), .B2(n480), .ZN(n3067) );
  OAI22_X1 U1656 ( .A1(n3679), .A2(n335), .B1(n74), .B2(n479), .ZN(n3068) );
  OAI22_X1 U1657 ( .A1(n3663), .A2(n336), .B1(n74), .B2(n478), .ZN(n3069) );
  OAI22_X1 U1658 ( .A1(n3647), .A2(n335), .B1(n74), .B2(n477), .ZN(n3070) );
  OAI22_X1 U1659 ( .A1(n3631), .A2(n336), .B1(n74), .B2(n476), .ZN(n3071) );
  OAI22_X1 U1660 ( .A1(n3615), .A2(n335), .B1(n74), .B2(n475), .ZN(n3072) );
  OAI22_X1 U1661 ( .A1(n3599), .A2(n336), .B1(n74), .B2(n474), .ZN(n3073) );
  OAI22_X1 U1662 ( .A1(n3583), .A2(n335), .B1(n74), .B2(n473), .ZN(n3074) );
  OAI22_X1 U1663 ( .A1(n3567), .A2(n336), .B1(n74), .B2(n472), .ZN(n3075) );
  OAI22_X1 U1664 ( .A1(n3551), .A2(n336), .B1(n74), .B2(n471), .ZN(n3076) );
  OAI22_X1 U1665 ( .A1(n3535), .A2(n336), .B1(n74), .B2(n470), .ZN(n3077) );
  OAI22_X1 U1666 ( .A1(n3519), .A2(n336), .B1(n74), .B2(n469), .ZN(n3078) );
  OAI22_X1 U1667 ( .A1(n3503), .A2(n336), .B1(n74), .B2(n468), .ZN(n3079) );
  OAI22_X1 U1668 ( .A1(n3487), .A2(n336), .B1(n74), .B2(n467), .ZN(n3080) );
  OAI22_X1 U1669 ( .A1(n3471), .A2(n336), .B1(n74), .B2(n466), .ZN(n3081) );
  OAI22_X1 U1670 ( .A1(n3455), .A2(n336), .B1(n74), .B2(n465), .ZN(n3082) );
  OAI22_X1 U1671 ( .A1(n3439), .A2(n336), .B1(n74), .B2(n464), .ZN(n3083) );
  OAI22_X1 U1672 ( .A1(n3423), .A2(n336), .B1(n74), .B2(n463), .ZN(n3084) );
  OAI22_X1 U1673 ( .A1(n3407), .A2(n336), .B1(n74), .B2(n462), .ZN(n3085) );
  OAI22_X1 U1674 ( .A1(n3391), .A2(n336), .B1(n74), .B2(n461), .ZN(n3086) );
  OAI22_X1 U1675 ( .A1(n3375), .A2(n335), .B1(n74), .B2(n460), .ZN(n3087) );
  OAI22_X1 U1676 ( .A1(n3359), .A2(n335), .B1(n74), .B2(n459), .ZN(n3088) );
  OAI22_X1 U1677 ( .A1(n3343), .A2(n335), .B1(n74), .B2(n458), .ZN(n3089) );
  OAI22_X1 U1678 ( .A1(n3327), .A2(n335), .B1(n74), .B2(n457), .ZN(n3090) );
  OAI22_X1 U1679 ( .A1(n3311), .A2(n335), .B1(n74), .B2(n456), .ZN(n3091) );
  OAI22_X1 U1680 ( .A1(n3295), .A2(n335), .B1(n74), .B2(n455), .ZN(n3092) );
  OAI22_X1 U1681 ( .A1(n2361), .A2(n335), .B1(n74), .B2(n454), .ZN(n3093) );
  OAI22_X1 U1682 ( .A1(n1058), .A2(n335), .B1(n74), .B2(n453), .ZN(n3094) );
  OAI22_X1 U1683 ( .A1(n1042), .A2(n335), .B1(n74), .B2(n452), .ZN(n3095) );
  OAI22_X1 U1684 ( .A1(n1026), .A2(n335), .B1(n74), .B2(n451), .ZN(n3096) );
  OAI22_X1 U1685 ( .A1(n1010), .A2(n335), .B1(n74), .B2(n450), .ZN(n3097) );
  OAI22_X1 U1686 ( .A1(n994), .A2(n335), .B1(n74), .B2(n449), .ZN(n3098) );
  OAI22_X1 U1687 ( .A1(n3695), .A2(n163), .B1(n75), .B2(n320), .ZN(n3099) );
  OAI22_X1 U1688 ( .A1(n3679), .A2(n162), .B1(n75), .B2(n319), .ZN(n3100) );
  OAI22_X1 U1689 ( .A1(n3663), .A2(n163), .B1(n75), .B2(n318), .ZN(n3101) );
  OAI22_X1 U1690 ( .A1(n3647), .A2(n162), .B1(n75), .B2(n317), .ZN(n3102) );
  OAI22_X1 U1691 ( .A1(n3631), .A2(n163), .B1(n75), .B2(n316), .ZN(n3103) );
  OAI22_X1 U1692 ( .A1(n3615), .A2(n162), .B1(n75), .B2(n315), .ZN(n3104) );
  OAI22_X1 U1693 ( .A1(n3599), .A2(n163), .B1(n75), .B2(n314), .ZN(n3105) );
  OAI22_X1 U1694 ( .A1(n3583), .A2(n162), .B1(n75), .B2(n313), .ZN(n3106) );
  OAI22_X1 U1695 ( .A1(n3567), .A2(n163), .B1(n75), .B2(n312), .ZN(n3107) );
  OAI22_X1 U1696 ( .A1(n3551), .A2(n163), .B1(n75), .B2(n311), .ZN(n3108) );
  OAI22_X1 U1697 ( .A1(n3535), .A2(n163), .B1(n75), .B2(n310), .ZN(n3109) );
  OAI22_X1 U1698 ( .A1(n3519), .A2(n163), .B1(n75), .B2(n309), .ZN(n3110) );
  OAI22_X1 U1699 ( .A1(n3503), .A2(n163), .B1(n75), .B2(n308), .ZN(n3111) );
  OAI22_X1 U1700 ( .A1(n3487), .A2(n163), .B1(n75), .B2(n307), .ZN(n3112) );
  OAI22_X1 U1701 ( .A1(n3471), .A2(n163), .B1(n75), .B2(n306), .ZN(n3113) );
  OAI22_X1 U1702 ( .A1(n3455), .A2(n163), .B1(n75), .B2(n305), .ZN(n3114) );
  OAI22_X1 U1703 ( .A1(n3439), .A2(n163), .B1(n75), .B2(n304), .ZN(n3115) );
  OAI22_X1 U1704 ( .A1(n3423), .A2(n163), .B1(n75), .B2(n303), .ZN(n3116) );
  OAI22_X1 U1705 ( .A1(n3407), .A2(n163), .B1(n75), .B2(n302), .ZN(n3117) );
  OAI22_X1 U1706 ( .A1(n3391), .A2(n163), .B1(n75), .B2(n301), .ZN(n3118) );
  OAI22_X1 U1707 ( .A1(n3375), .A2(n162), .B1(n75), .B2(n300), .ZN(n3119) );
  OAI22_X1 U1708 ( .A1(n3359), .A2(n162), .B1(n75), .B2(n299), .ZN(n3120) );
  OAI22_X1 U1709 ( .A1(n3343), .A2(n162), .B1(n75), .B2(n298), .ZN(n3121) );
  OAI22_X1 U1710 ( .A1(n3327), .A2(n162), .B1(n75), .B2(n297), .ZN(n3122) );
  OAI22_X1 U1711 ( .A1(n3311), .A2(n162), .B1(n75), .B2(n296), .ZN(n3123) );
  OAI22_X1 U1712 ( .A1(n3295), .A2(n162), .B1(n75), .B2(n295), .ZN(n3124) );
  OAI22_X1 U1713 ( .A1(n2361), .A2(n162), .B1(n75), .B2(n294), .ZN(n3125) );
  OAI22_X1 U1714 ( .A1(n1058), .A2(n162), .B1(n75), .B2(n293), .ZN(n3126) );
  OAI22_X1 U1715 ( .A1(n1042), .A2(n162), .B1(n75), .B2(n292), .ZN(n3127) );
  OAI22_X1 U1716 ( .A1(n1026), .A2(n162), .B1(n75), .B2(n291), .ZN(n3128) );
  OAI22_X1 U1717 ( .A1(n1010), .A2(n162), .B1(n75), .B2(n290), .ZN(n3129) );
  OAI22_X1 U1718 ( .A1(n994), .A2(n162), .B1(n75), .B2(n289), .ZN(n3130) );
  OAI22_X1 U1719 ( .A1(n3695), .A2(n154), .B1(n68), .B2(n288), .ZN(n3131) );
  OAI22_X1 U1720 ( .A1(n3679), .A2(n153), .B1(n68), .B2(n287), .ZN(n3132) );
  OAI22_X1 U1721 ( .A1(n3663), .A2(n154), .B1(n68), .B2(n286), .ZN(n3133) );
  OAI22_X1 U1722 ( .A1(n3647), .A2(n153), .B1(n68), .B2(n285), .ZN(n3134) );
  OAI22_X1 U1723 ( .A1(n3631), .A2(n154), .B1(n68), .B2(n284), .ZN(n3135) );
  OAI22_X1 U1724 ( .A1(n3615), .A2(n153), .B1(n68), .B2(n283), .ZN(n3136) );
  OAI22_X1 U1725 ( .A1(n3599), .A2(n154), .B1(n68), .B2(n282), .ZN(n3137) );
  OAI22_X1 U1726 ( .A1(n3583), .A2(n153), .B1(n68), .B2(n281), .ZN(n3138) );
  OAI22_X1 U1727 ( .A1(n3567), .A2(n154), .B1(n68), .B2(n280), .ZN(n3139) );
  OAI22_X1 U1728 ( .A1(n3551), .A2(n154), .B1(n68), .B2(n279), .ZN(n3140) );
  OAI22_X1 U1729 ( .A1(n3535), .A2(n154), .B1(n68), .B2(n278), .ZN(n3141) );
  OAI22_X1 U1730 ( .A1(n3519), .A2(n154), .B1(n68), .B2(n277), .ZN(n3142) );
  OAI22_X1 U1731 ( .A1(n3503), .A2(n154), .B1(n68), .B2(n276), .ZN(n3143) );
  OAI22_X1 U1732 ( .A1(n3487), .A2(n154), .B1(n68), .B2(n275), .ZN(n3144) );
  OAI22_X1 U1733 ( .A1(n3471), .A2(n154), .B1(n68), .B2(n274), .ZN(n3145) );
  OAI22_X1 U1734 ( .A1(n3455), .A2(n154), .B1(n68), .B2(n273), .ZN(n3146) );
  OAI22_X1 U1735 ( .A1(n3439), .A2(n154), .B1(n68), .B2(n272), .ZN(n3147) );
  OAI22_X1 U1736 ( .A1(n3423), .A2(n154), .B1(n68), .B2(n271), .ZN(n3148) );
  OAI22_X1 U1737 ( .A1(n3407), .A2(n154), .B1(n68), .B2(n270), .ZN(n3149) );
  OAI22_X1 U1738 ( .A1(n3391), .A2(n154), .B1(n68), .B2(n269), .ZN(n3150) );
  OAI22_X1 U1739 ( .A1(n3375), .A2(n153), .B1(n68), .B2(n268), .ZN(n3151) );
  OAI22_X1 U1740 ( .A1(n3359), .A2(n153), .B1(n68), .B2(n267), .ZN(n3152) );
  OAI22_X1 U1741 ( .A1(n3343), .A2(n153), .B1(n68), .B2(n266), .ZN(n3153) );
  OAI22_X1 U1742 ( .A1(n3327), .A2(n153), .B1(n68), .B2(n265), .ZN(n3154) );
  OAI22_X1 U1743 ( .A1(n3311), .A2(n153), .B1(n68), .B2(n264), .ZN(n3155) );
  OAI22_X1 U1744 ( .A1(n3295), .A2(n153), .B1(n68), .B2(n263), .ZN(n3156) );
  OAI22_X1 U1745 ( .A1(n2361), .A2(n153), .B1(n68), .B2(n262), .ZN(n3157) );
  OAI22_X1 U1746 ( .A1(n1058), .A2(n153), .B1(n68), .B2(n261), .ZN(n3158) );
  OAI22_X1 U1747 ( .A1(n1042), .A2(n153), .B1(n68), .B2(n260), .ZN(n3159) );
  OAI22_X1 U1748 ( .A1(n1026), .A2(n153), .B1(n68), .B2(n259), .ZN(n3160) );
  OAI22_X1 U1749 ( .A1(n1010), .A2(n153), .B1(n68), .B2(n258), .ZN(n3161) );
  OAI22_X1 U1750 ( .A1(n994), .A2(n153), .B1(n68), .B2(n257), .ZN(n3162) );
  OAI22_X1 U1751 ( .A1(n3695), .A2(n145), .B1(n67), .B2(n256), .ZN(n3163) );
  OAI22_X1 U1752 ( .A1(n3679), .A2(n144), .B1(n67), .B2(n255), .ZN(n3164) );
  OAI22_X1 U1753 ( .A1(n3663), .A2(n145), .B1(n67), .B2(n254), .ZN(n3165) );
  OAI22_X1 U1754 ( .A1(n3647), .A2(n144), .B1(n67), .B2(n253), .ZN(n3166) );
  OAI22_X1 U1755 ( .A1(n3631), .A2(n145), .B1(n67), .B2(n252), .ZN(n3167) );
  OAI22_X1 U1756 ( .A1(n3615), .A2(n144), .B1(n67), .B2(n251), .ZN(n3168) );
  OAI22_X1 U1757 ( .A1(n3599), .A2(n145), .B1(n67), .B2(n250), .ZN(n3169) );
  OAI22_X1 U1758 ( .A1(n3583), .A2(n144), .B1(n67), .B2(n249), .ZN(n3170) );
  OAI22_X1 U1759 ( .A1(n3567), .A2(n145), .B1(n67), .B2(n248), .ZN(n3171) );
  OAI22_X1 U1760 ( .A1(n3551), .A2(n145), .B1(n67), .B2(n247), .ZN(n3172) );
  OAI22_X1 U1761 ( .A1(n3535), .A2(n145), .B1(n67), .B2(n246), .ZN(n3173) );
  OAI22_X1 U1762 ( .A1(n3519), .A2(n145), .B1(n67), .B2(n245), .ZN(n3174) );
  OAI22_X1 U1763 ( .A1(n3503), .A2(n145), .B1(n67), .B2(n244), .ZN(n3175) );
  OAI22_X1 U1764 ( .A1(n3487), .A2(n145), .B1(n67), .B2(n243), .ZN(n3176) );
  OAI22_X1 U1765 ( .A1(n3471), .A2(n145), .B1(n67), .B2(n242), .ZN(n3177) );
  OAI22_X1 U1766 ( .A1(n3455), .A2(n145), .B1(n67), .B2(n241), .ZN(n3178) );
  OAI22_X1 U1767 ( .A1(n3439), .A2(n145), .B1(n67), .B2(n240), .ZN(n3179) );
  OAI22_X1 U1768 ( .A1(n3423), .A2(n145), .B1(n67), .B2(n239), .ZN(n3180) );
  OAI22_X1 U1769 ( .A1(n3407), .A2(n145), .B1(n67), .B2(n238), .ZN(n3181) );
  OAI22_X1 U1770 ( .A1(n3391), .A2(n145), .B1(n67), .B2(n237), .ZN(n3182) );
  OAI22_X1 U1771 ( .A1(n3375), .A2(n144), .B1(n67), .B2(n236), .ZN(n3183) );
  OAI22_X1 U1772 ( .A1(n3359), .A2(n144), .B1(n67), .B2(n235), .ZN(n3184) );
  OAI22_X1 U1773 ( .A1(n3343), .A2(n144), .B1(n67), .B2(n234), .ZN(n3185) );
  OAI22_X1 U1774 ( .A1(n3327), .A2(n144), .B1(n67), .B2(n233), .ZN(n3186) );
  OAI22_X1 U1775 ( .A1(n3311), .A2(n144), .B1(n67), .B2(n232), .ZN(n3187) );
  OAI22_X1 U1776 ( .A1(n3295), .A2(n144), .B1(n67), .B2(n231), .ZN(n3188) );
  OAI22_X1 U1777 ( .A1(n2361), .A2(n144), .B1(n67), .B2(n230), .ZN(n3189) );
  OAI22_X1 U1778 ( .A1(n1058), .A2(n144), .B1(n67), .B2(n229), .ZN(n3190) );
  OAI22_X1 U1779 ( .A1(n1042), .A2(n144), .B1(n67), .B2(n228), .ZN(n3191) );
  OAI22_X1 U1780 ( .A1(n1026), .A2(n144), .B1(n67), .B2(n227), .ZN(n3192) );
  OAI22_X1 U1781 ( .A1(n1010), .A2(n144), .B1(n67), .B2(n226), .ZN(n3193) );
  OAI22_X1 U1782 ( .A1(n994), .A2(n144), .B1(n67), .B2(n225), .ZN(n3194) );
  OAI22_X1 U1783 ( .A1(n3695), .A2(n136), .B1(n76), .B2(n224), .ZN(n3195) );
  OAI22_X1 U1784 ( .A1(n3679), .A2(n135), .B1(n76), .B2(n223), .ZN(n3196) );
  OAI22_X1 U1785 ( .A1(n3663), .A2(n136), .B1(n76), .B2(n222), .ZN(n3197) );
  OAI22_X1 U1786 ( .A1(n3647), .A2(n135), .B1(n76), .B2(n221), .ZN(n3198) );
  OAI22_X1 U1787 ( .A1(n3631), .A2(n136), .B1(n76), .B2(n220), .ZN(n3199) );
  OAI22_X1 U1788 ( .A1(n3615), .A2(n135), .B1(n76), .B2(n219), .ZN(n3200) );
  OAI22_X1 U1789 ( .A1(n3599), .A2(n136), .B1(n76), .B2(n218), .ZN(n3201) );
  OAI22_X1 U1790 ( .A1(n3583), .A2(n135), .B1(n76), .B2(n217), .ZN(n3202) );
  OAI22_X1 U1791 ( .A1(n3567), .A2(n136), .B1(n76), .B2(n216), .ZN(n3203) );
  OAI22_X1 U1792 ( .A1(n3551), .A2(n136), .B1(n76), .B2(n215), .ZN(n3204) );
  OAI22_X1 U1793 ( .A1(n3535), .A2(n136), .B1(n76), .B2(n214), .ZN(n3205) );
  OAI22_X1 U1794 ( .A1(n3519), .A2(n136), .B1(n76), .B2(n213), .ZN(n3206) );
  OAI22_X1 U1795 ( .A1(n3503), .A2(n136), .B1(n76), .B2(n212), .ZN(n3207) );
  OAI22_X1 U1796 ( .A1(n3487), .A2(n136), .B1(n76), .B2(n211), .ZN(n3208) );
  OAI22_X1 U1797 ( .A1(n3471), .A2(n136), .B1(n76), .B2(n210), .ZN(n3209) );
  OAI22_X1 U1798 ( .A1(n3455), .A2(n136), .B1(n76), .B2(n209), .ZN(n3210) );
  OAI22_X1 U1799 ( .A1(n3439), .A2(n136), .B1(n76), .B2(n208), .ZN(n3211) );
  OAI22_X1 U1800 ( .A1(n3423), .A2(n136), .B1(n76), .B2(n207), .ZN(n3212) );
  OAI22_X1 U1801 ( .A1(n3407), .A2(n136), .B1(n76), .B2(n206), .ZN(n3213) );
  OAI22_X1 U1802 ( .A1(n3391), .A2(n136), .B1(n76), .B2(n205), .ZN(n3214) );
  OAI22_X1 U1803 ( .A1(n3375), .A2(n135), .B1(n76), .B2(n204), .ZN(n3215) );
  OAI22_X1 U1804 ( .A1(n3359), .A2(n135), .B1(n76), .B2(n203), .ZN(n3216) );
  OAI22_X1 U1805 ( .A1(n3343), .A2(n135), .B1(n76), .B2(n202), .ZN(n3217) );
  OAI22_X1 U1806 ( .A1(n3327), .A2(n135), .B1(n76), .B2(n201), .ZN(n3218) );
  OAI22_X1 U1807 ( .A1(n3311), .A2(n135), .B1(n76), .B2(n200), .ZN(n3219) );
  OAI22_X1 U1808 ( .A1(n3295), .A2(n135), .B1(n76), .B2(n199), .ZN(n3220) );
  OAI22_X1 U1809 ( .A1(n2361), .A2(n135), .B1(n76), .B2(n198), .ZN(n3221) );
  OAI22_X1 U1810 ( .A1(n1058), .A2(n135), .B1(n76), .B2(n197), .ZN(n3222) );
  OAI22_X1 U1811 ( .A1(n1042), .A2(n135), .B1(n76), .B2(n196), .ZN(n3223) );
  OAI22_X1 U1812 ( .A1(n1026), .A2(n135), .B1(n76), .B2(n195), .ZN(n3224) );
  OAI22_X1 U1813 ( .A1(n1010), .A2(n135), .B1(n76), .B2(n194), .ZN(n3225) );
  OAI22_X1 U1814 ( .A1(n994), .A2(n135), .B1(n76), .B2(n193), .ZN(n3226) );
  OAI22_X1 U1815 ( .A1(n3695), .A2(n91), .B1(n77), .B2(n64), .ZN(n3227) );
  OAI22_X1 U1816 ( .A1(n3679), .A2(n90), .B1(n77), .B2(n63), .ZN(n3228) );
  OAI22_X1 U1817 ( .A1(n3663), .A2(n91), .B1(n77), .B2(n62), .ZN(n3229) );
  OAI22_X1 U1818 ( .A1(n3647), .A2(n90), .B1(n77), .B2(n61), .ZN(n3230) );
  OAI22_X1 U1819 ( .A1(n3631), .A2(n91), .B1(n77), .B2(n60), .ZN(n3231) );
  OAI22_X1 U1820 ( .A1(n3615), .A2(n90), .B1(n77), .B2(n59), .ZN(n3232) );
  OAI22_X1 U1821 ( .A1(n3599), .A2(n91), .B1(n77), .B2(n58), .ZN(n3233) );
  OAI22_X1 U1822 ( .A1(n3583), .A2(n90), .B1(n77), .B2(n57), .ZN(n3234) );
  OAI22_X1 U1823 ( .A1(n3567), .A2(n91), .B1(n77), .B2(n56), .ZN(n3235) );
  OAI22_X1 U1824 ( .A1(n3551), .A2(n91), .B1(n77), .B2(n55), .ZN(n3236) );
  OAI22_X1 U1825 ( .A1(n3535), .A2(n91), .B1(n77), .B2(n54), .ZN(n3237) );
  OAI22_X1 U1826 ( .A1(n3519), .A2(n91), .B1(n77), .B2(n53), .ZN(n3238) );
  OAI22_X1 U1827 ( .A1(n3503), .A2(n91), .B1(n77), .B2(n52), .ZN(n3239) );
  OAI22_X1 U1828 ( .A1(n3487), .A2(n91), .B1(n77), .B2(n51), .ZN(n3240) );
  OAI22_X1 U1829 ( .A1(n3471), .A2(n91), .B1(n77), .B2(n50), .ZN(n3241) );
  OAI22_X1 U1830 ( .A1(n3455), .A2(n91), .B1(n77), .B2(n49), .ZN(n3242) );
  OAI22_X1 U1831 ( .A1(n3439), .A2(n91), .B1(n77), .B2(n48), .ZN(n3243) );
  OAI22_X1 U1832 ( .A1(n3423), .A2(n91), .B1(n77), .B2(n47), .ZN(n3244) );
  OAI22_X1 U1833 ( .A1(n3407), .A2(n91), .B1(n77), .B2(n46), .ZN(n3245) );
  OAI22_X1 U1834 ( .A1(n3391), .A2(n91), .B1(n77), .B2(n45), .ZN(n3246) );
  OAI22_X1 U1835 ( .A1(n3375), .A2(n90), .B1(n77), .B2(n44), .ZN(n3247) );
  OAI22_X1 U1836 ( .A1(n3359), .A2(n90), .B1(n77), .B2(n43), .ZN(n3248) );
  OAI22_X1 U1837 ( .A1(n3343), .A2(n90), .B1(n77), .B2(n42), .ZN(n3249) );
  OAI22_X1 U1838 ( .A1(n3327), .A2(n90), .B1(n77), .B2(n41), .ZN(n3250) );
  OAI22_X1 U1839 ( .A1(n3311), .A2(n90), .B1(n77), .B2(n40), .ZN(n3251) );
  OAI22_X1 U1840 ( .A1(n3295), .A2(n90), .B1(n77), .B2(n39), .ZN(n3252) );
  OAI22_X1 U1841 ( .A1(n2361), .A2(n90), .B1(n77), .B2(n38), .ZN(n3253) );
  OAI22_X1 U1842 ( .A1(n1058), .A2(n90), .B1(n77), .B2(n37), .ZN(n3254) );
  OAI22_X1 U1843 ( .A1(n1042), .A2(n90), .B1(n77), .B2(n36), .ZN(n3255) );
  OAI22_X1 U1844 ( .A1(n1026), .A2(n90), .B1(n77), .B2(n35), .ZN(n3256) );
  OAI22_X1 U1845 ( .A1(n1010), .A2(n90), .B1(n77), .B2(n34), .ZN(n3257) );
  OAI22_X1 U1846 ( .A1(n994), .A2(n90), .B1(n77), .B2(n33), .ZN(n3258) );
  OAI22_X1 U1847 ( .A1(n3695), .A2(n82), .B1(n80), .B2(n32), .ZN(n3259) );
  OAI22_X1 U1848 ( .A1(n3679), .A2(n81), .B1(n80), .B2(n31), .ZN(n3260) );
  OAI22_X1 U1849 ( .A1(n3663), .A2(n82), .B1(n80), .B2(n30), .ZN(n3261) );
  OAI22_X1 U1850 ( .A1(n3647), .A2(n81), .B1(n80), .B2(n29), .ZN(n3262) );
  OAI22_X1 U1851 ( .A1(n3631), .A2(n82), .B1(n80), .B2(n28), .ZN(n3263) );
  OAI22_X1 U1852 ( .A1(n3615), .A2(n81), .B1(n80), .B2(n27), .ZN(n3264) );
  OAI22_X1 U1853 ( .A1(n3599), .A2(n82), .B1(n80), .B2(n26), .ZN(n3265) );
  OAI22_X1 U1854 ( .A1(n3583), .A2(n81), .B1(n80), .B2(n25), .ZN(n3266) );
  OAI22_X1 U1855 ( .A1(n3567), .A2(n82), .B1(n80), .B2(n24), .ZN(n3267) );
  OAI22_X1 U1856 ( .A1(n3551), .A2(n82), .B1(n80), .B2(n23), .ZN(n3268) );
  OAI22_X1 U1857 ( .A1(n3535), .A2(n82), .B1(n80), .B2(n22), .ZN(n3269) );
  OAI22_X1 U1858 ( .A1(n3519), .A2(n82), .B1(n80), .B2(n21), .ZN(n3270) );
  OAI22_X1 U1859 ( .A1(n3503), .A2(n82), .B1(n80), .B2(n20), .ZN(n3271) );
  OAI22_X1 U1860 ( .A1(n3487), .A2(n82), .B1(n80), .B2(n19), .ZN(n3272) );
  OAI22_X1 U1861 ( .A1(n3471), .A2(n82), .B1(n80), .B2(n18), .ZN(n3273) );
  OAI22_X1 U1862 ( .A1(n3455), .A2(n82), .B1(n80), .B2(n17), .ZN(n3274) );
  OAI22_X1 U1863 ( .A1(n3439), .A2(n82), .B1(n80), .B2(n16), .ZN(n3275) );
  OAI22_X1 U1864 ( .A1(n3423), .A2(n82), .B1(n80), .B2(n15), .ZN(n3276) );
  OAI22_X1 U1865 ( .A1(n3407), .A2(n82), .B1(n80), .B2(n14), .ZN(n3277) );
  OAI22_X1 U1866 ( .A1(n3391), .A2(n82), .B1(n80), .B2(n13), .ZN(n3278) );
  OAI22_X1 U1867 ( .A1(n3375), .A2(n81), .B1(n80), .B2(n12), .ZN(n3279) );
  OAI22_X1 U1868 ( .A1(n3359), .A2(n81), .B1(n80), .B2(n11), .ZN(n3280) );
  OAI22_X1 U1869 ( .A1(n3343), .A2(n81), .B1(n80), .B2(n10), .ZN(n3281) );
  OAI22_X1 U1870 ( .A1(n3327), .A2(n81), .B1(n80), .B2(n9), .ZN(n3282) );
  OAI22_X1 U1871 ( .A1(n3311), .A2(n81), .B1(n80), .B2(n8), .ZN(n3283) );
  OAI22_X1 U1872 ( .A1(n3295), .A2(n81), .B1(n80), .B2(n7), .ZN(n3284) );
  OAI22_X1 U1873 ( .A1(n2361), .A2(n81), .B1(n80), .B2(n6), .ZN(n3285) );
  OAI22_X1 U1874 ( .A1(n1058), .A2(n81), .B1(n80), .B2(n5), .ZN(n3286) );
  OAI22_X1 U1875 ( .A1(n1042), .A2(n81), .B1(n80), .B2(n4), .ZN(n3287) );
  OAI22_X1 U1876 ( .A1(n1026), .A2(n81), .B1(n80), .B2(n3), .ZN(n3288) );
  OAI22_X1 U1877 ( .A1(n1010), .A2(n81), .B1(n80), .B2(n2), .ZN(n3289) );
  OAI22_X1 U1878 ( .A1(n994), .A2(n81), .B1(n80), .B2(n1), .ZN(n3290) );
  NOR2_X1 U1879 ( .A1(wa[2]), .A2(wa[3]), .ZN(n2430) );
  NOR2_X1 U1880 ( .A1(n3711), .A2(wa[2]), .ZN(n2571) );
  NOR2_X1 U1881 ( .A1(n3712), .A2(wa[3]), .ZN(n2359) );
  AOI221_X1 U1882 ( .B1(x9_s1_w[0]), .B2(n1113), .C1(x8_s0_w[0]), .C2(n1114), 
        .A(n1658), .ZN(n1628) );
  AOI221_X1 U1883 ( .B1(x15_a5_w[0]), .B2(n1108), .C1(x14_a4_w[0]), .C2(n1109), 
        .A(n1657), .ZN(n1629) );
  AOI211_X1 U1884 ( .C1(x1_ra_w[0]), .C2(n1098), .A(n1650), .B(n1651), .ZN(
        n1630) );
  AOI221_X1 U1885 ( .B1(x9_s1_w[1]), .B2(n1113), .C1(x8_s0_w[1]), .C2(n1114), 
        .A(n1457), .ZN(n1441) );
  AOI221_X1 U1886 ( .B1(x15_a5_w[1]), .B2(n1108), .C1(x14_a4_w[1]), .C2(n1109), 
        .A(n1456), .ZN(n1442) );
  AOI211_X1 U1887 ( .C1(x1_ra_w[1]), .C2(n1098), .A(n1453), .B(n1454), .ZN(
        n1443) );
  AOI221_X1 U1888 ( .B1(x9_s1_w[2]), .B2(n1113), .C1(x8_s0_w[2]), .C2(n1114), 
        .A(n1270), .ZN(n1254) );
  AOI221_X1 U1889 ( .B1(x15_a5_w[2]), .B2(n1108), .C1(x14_a4_w[2]), .C2(n1109), 
        .A(n1269), .ZN(n1255) );
  AOI211_X1 U1890 ( .C1(x1_ra_w[2]), .C2(n1098), .A(n1266), .B(n1267), .ZN(
        n1256) );
  AOI221_X1 U1891 ( .B1(x9_s1_w[3]), .B2(n1113), .C1(x8_s0_w[3]), .C2(n1114), 
        .A(n1219), .ZN(n1203) );
  AOI221_X1 U1892 ( .B1(x15_a5_w[3]), .B2(n1108), .C1(x14_a4_w[3]), .C2(n1109), 
        .A(n1218), .ZN(n1204) );
  AOI211_X1 U1893 ( .C1(x1_ra_w[3]), .C2(n1098), .A(n1215), .B(n1216), .ZN(
        n1205) );
  AOI221_X1 U1894 ( .B1(x9_s1_w[4]), .B2(n1113), .C1(x8_s0_w[4]), .C2(n1114), 
        .A(n1202), .ZN(n1186) );
  AOI221_X1 U1895 ( .B1(x15_a5_w[4]), .B2(n1108), .C1(x14_a4_w[4]), .C2(n1109), 
        .A(n1201), .ZN(n1187) );
  AOI211_X1 U1896 ( .C1(x1_ra_w[4]), .C2(n1098), .A(n1198), .B(n1199), .ZN(
        n1188) );
  AOI221_X1 U1897 ( .B1(x9_s1_w[5]), .B2(n1113), .C1(x8_s0_w[5]), .C2(n1114), 
        .A(n1185), .ZN(n1169) );
  AOI221_X1 U1898 ( .B1(x15_a5_w[5]), .B2(n1108), .C1(x14_a4_w[5]), .C2(n1109), 
        .A(n1184), .ZN(n1170) );
  AOI211_X1 U1899 ( .C1(x1_ra_w[5]), .C2(n1098), .A(n1181), .B(n1182), .ZN(
        n1171) );
  AOI221_X1 U1900 ( .B1(x9_s1_w[6]), .B2(n1113), .C1(x8_s0_w[6]), .C2(n1114), 
        .A(n1168), .ZN(n1152) );
  AOI221_X1 U1901 ( .B1(x15_a5_w[6]), .B2(n1108), .C1(x14_a4_w[6]), .C2(n1109), 
        .A(n1167), .ZN(n1153) );
  AOI211_X1 U1902 ( .C1(x1_ra_w[6]), .C2(n1098), .A(n1164), .B(n1165), .ZN(
        n1154) );
  AOI221_X1 U1903 ( .B1(x9_s1_w[7]), .B2(n1113), .C1(x8_s0_w[7]), .C2(n1114), 
        .A(n1151), .ZN(n1135) );
  AOI221_X1 U1904 ( .B1(x15_a5_w[7]), .B2(n1108), .C1(x14_a4_w[7]), .C2(n1109), 
        .A(n1150), .ZN(n1136) );
  AOI211_X1 U1905 ( .C1(x1_ra_w[7]), .C2(n1098), .A(n1147), .B(n1148), .ZN(
        n1137) );
  AOI221_X1 U1906 ( .B1(x9_s1_w[8]), .B2(n1113), .C1(x8_s0_w[8]), .C2(n1114), 
        .A(n1134), .ZN(n1118) );
  AOI221_X1 U1907 ( .B1(x15_a5_w[8]), .B2(n1108), .C1(x14_a4_w[8]), .C2(n1109), 
        .A(n1133), .ZN(n1119) );
  AOI211_X1 U1908 ( .C1(x1_ra_w[8]), .C2(n1098), .A(n1130), .B(n1131), .ZN(
        n1120) );
  AOI221_X1 U1909 ( .B1(x9_s1_w[9]), .B2(n1113), .C1(x8_s0_w[9]), .C2(n1114), 
        .A(n1115), .ZN(n1070) );
  AOI221_X1 U1910 ( .B1(x15_a5_w[9]), .B2(n1108), .C1(x14_a4_w[9]), .C2(n1109), 
        .A(n1110), .ZN(n1071) );
  AOI211_X1 U1911 ( .C1(x1_ra_w[9]), .C2(n1098), .A(n1099), .B(n1100), .ZN(
        n1072) );
  AOI221_X1 U1912 ( .B1(x9_s1_w[10]), .B2(n1113), .C1(x8_s0_w[10]), .C2(n1114), 
        .A(n1627), .ZN(n1611) );
  AOI221_X1 U1913 ( .B1(x15_a5_w[10]), .B2(n1108), .C1(x14_a4_w[10]), .C2(
        n1109), .A(n1626), .ZN(n1612) );
  AOI211_X1 U1914 ( .C1(x1_ra_w[10]), .C2(n1098), .A(n1623), .B(n1624), .ZN(
        n1613) );
  AOI221_X1 U1915 ( .B1(x9_s1_w[11]), .B2(n1113), .C1(x8_s0_w[11]), .C2(n1114), 
        .A(n1610), .ZN(n1594) );
  AOI221_X1 U1916 ( .B1(x15_a5_w[11]), .B2(n1108), .C1(x14_a4_w[11]), .C2(
        n1109), .A(n1609), .ZN(n1595) );
  AOI211_X1 U1917 ( .C1(x1_ra_w[11]), .C2(n1098), .A(n1606), .B(n1607), .ZN(
        n1596) );
  AOI221_X1 U1918 ( .B1(x9_s1_w[12]), .B2(n1113), .C1(x8_s0_w[12]), .C2(n1114), 
        .A(n1593), .ZN(n1577) );
  AOI221_X1 U1919 ( .B1(x15_a5_w[12]), .B2(n1108), .C1(x14_a4_w[12]), .C2(
        n1109), .A(n1592), .ZN(n1578) );
  AOI211_X1 U1920 ( .C1(x1_ra_w[12]), .C2(n1098), .A(n1589), .B(n1590), .ZN(
        n1579) );
  AOI221_X1 U1921 ( .B1(x9_s1_w[13]), .B2(n1113), .C1(x8_s0_w[13]), .C2(n1114), 
        .A(n1576), .ZN(n1560) );
  AOI221_X1 U1922 ( .B1(x15_a5_w[13]), .B2(n1108), .C1(x14_a4_w[13]), .C2(
        n1109), .A(n1575), .ZN(n1561) );
  AOI211_X1 U1923 ( .C1(x1_ra_w[13]), .C2(n1098), .A(n1572), .B(n1573), .ZN(
        n1562) );
  AOI221_X1 U1924 ( .B1(x9_s1_w[14]), .B2(n1113), .C1(x8_s0_w[14]), .C2(n1114), 
        .A(n1559), .ZN(n1543) );
  AOI221_X1 U1925 ( .B1(x15_a5_w[14]), .B2(n1108), .C1(x14_a4_w[14]), .C2(
        n1109), .A(n1558), .ZN(n1544) );
  AOI211_X1 U1926 ( .C1(x1_ra_w[14]), .C2(n1098), .A(n1555), .B(n1556), .ZN(
        n1545) );
  AOI221_X1 U1927 ( .B1(x9_s1_w[15]), .B2(n1113), .C1(x8_s0_w[15]), .C2(n1114), 
        .A(n1542), .ZN(n1526) );
  AOI221_X1 U1928 ( .B1(x15_a5_w[15]), .B2(n1108), .C1(x14_a4_w[15]), .C2(
        n1109), .A(n1541), .ZN(n1527) );
  AOI211_X1 U1929 ( .C1(x1_ra_w[15]), .C2(n1098), .A(n1538), .B(n1539), .ZN(
        n1528) );
  AOI221_X1 U1930 ( .B1(x9_s1_w[16]), .B2(n1113), .C1(x8_s0_w[16]), .C2(n1114), 
        .A(n1525), .ZN(n1509) );
  AOI221_X1 U1931 ( .B1(x15_a5_w[16]), .B2(n1108), .C1(x14_a4_w[16]), .C2(
        n1109), .A(n1524), .ZN(n1510) );
  AOI211_X1 U1932 ( .C1(x1_ra_w[16]), .C2(n1098), .A(n1521), .B(n1522), .ZN(
        n1511) );
  AOI221_X1 U1933 ( .B1(x9_s1_w[17]), .B2(n1113), .C1(x8_s0_w[17]), .C2(n1114), 
        .A(n1508), .ZN(n1492) );
  AOI221_X1 U1934 ( .B1(x15_a5_w[17]), .B2(n1108), .C1(x14_a4_w[17]), .C2(
        n1109), .A(n1507), .ZN(n1493) );
  AOI211_X1 U1935 ( .C1(x1_ra_w[17]), .C2(n1098), .A(n1504), .B(n1505), .ZN(
        n1494) );
  AOI221_X1 U1936 ( .B1(x9_s1_w[18]), .B2(n1113), .C1(x8_s0_w[18]), .C2(n1114), 
        .A(n1491), .ZN(n1475) );
  AOI221_X1 U1937 ( .B1(x15_a5_w[18]), .B2(n1108), .C1(x14_a4_w[18]), .C2(
        n1109), .A(n1490), .ZN(n1476) );
  AOI211_X1 U1938 ( .C1(x1_ra_w[18]), .C2(n1098), .A(n1487), .B(n1488), .ZN(
        n1477) );
  AOI221_X1 U1939 ( .B1(x9_s1_w[19]), .B2(n1113), .C1(x8_s0_w[19]), .C2(n1114), 
        .A(n1474), .ZN(n1458) );
  AOI221_X1 U1940 ( .B1(x15_a5_w[19]), .B2(n1108), .C1(x14_a4_w[19]), .C2(
        n1109), .A(n1473), .ZN(n1459) );
  AOI211_X1 U1941 ( .C1(x1_ra_w[19]), .C2(n1098), .A(n1470), .B(n1471), .ZN(
        n1460) );
  AOI221_X1 U1942 ( .B1(x9_s1_w[20]), .B2(n1113), .C1(x8_s0_w[20]), .C2(n1114), 
        .A(n1440), .ZN(n1424) );
  AOI221_X1 U1943 ( .B1(x15_a5_w[20]), .B2(n1108), .C1(x14_a4_w[20]), .C2(
        n1109), .A(n1439), .ZN(n1425) );
  AOI211_X1 U1944 ( .C1(x1_ra_w[20]), .C2(n1098), .A(n1436), .B(n1437), .ZN(
        n1426) );
  AOI221_X1 U1945 ( .B1(x9_s1_w[21]), .B2(n1113), .C1(x8_s0_w[21]), .C2(n1114), 
        .A(n1423), .ZN(n1407) );
  AOI221_X1 U1946 ( .B1(x15_a5_w[21]), .B2(n1108), .C1(x14_a4_w[21]), .C2(
        n1109), .A(n1422), .ZN(n1408) );
  AOI211_X1 U1947 ( .C1(x1_ra_w[21]), .C2(n1098), .A(n1419), .B(n1420), .ZN(
        n1409) );
  AOI221_X1 U1948 ( .B1(x9_s1_w[22]), .B2(n1113), .C1(x8_s0_w[22]), .C2(n1114), 
        .A(n1406), .ZN(n1390) );
  AOI221_X1 U1949 ( .B1(x15_a5_w[22]), .B2(n1108), .C1(x14_a4_w[22]), .C2(
        n1109), .A(n1405), .ZN(n1391) );
  AOI211_X1 U1950 ( .C1(x1_ra_w[22]), .C2(n1098), .A(n1402), .B(n1403), .ZN(
        n1392) );
  AOI221_X1 U1951 ( .B1(x9_s1_w[23]), .B2(n1113), .C1(x8_s0_w[23]), .C2(n1114), 
        .A(n1389), .ZN(n1373) );
  AOI221_X1 U1952 ( .B1(x15_a5_w[23]), .B2(n1108), .C1(x14_a4_w[23]), .C2(
        n1109), .A(n1388), .ZN(n1374) );
  AOI211_X1 U1953 ( .C1(x1_ra_w[23]), .C2(n1098), .A(n1385), .B(n1386), .ZN(
        n1375) );
  AOI221_X1 U1954 ( .B1(x9_s1_w[24]), .B2(n1113), .C1(x8_s0_w[24]), .C2(n1114), 
        .A(n1372), .ZN(n1356) );
  AOI221_X1 U1955 ( .B1(x15_a5_w[24]), .B2(n1108), .C1(x14_a4_w[24]), .C2(
        n1109), .A(n1371), .ZN(n1357) );
  AOI211_X1 U1956 ( .C1(x1_ra_w[24]), .C2(n1098), .A(n1368), .B(n1369), .ZN(
        n1358) );
  AOI221_X1 U1957 ( .B1(x9_s1_w[25]), .B2(n1113), .C1(x8_s0_w[25]), .C2(n1114), 
        .A(n1355), .ZN(n1339) );
  AOI221_X1 U1958 ( .B1(x15_a5_w[25]), .B2(n1108), .C1(x14_a4_w[25]), .C2(
        n1109), .A(n1354), .ZN(n1340) );
  AOI211_X1 U1959 ( .C1(x1_ra_w[25]), .C2(n1098), .A(n1351), .B(n1352), .ZN(
        n1341) );
  AOI221_X1 U1960 ( .B1(x9_s1_w[26]), .B2(n1113), .C1(x8_s0_w[26]), .C2(n1114), 
        .A(n1338), .ZN(n1322) );
  AOI221_X1 U1961 ( .B1(x15_a5_w[26]), .B2(n1108), .C1(x14_a4_w[26]), .C2(
        n1109), .A(n1337), .ZN(n1323) );
  AOI211_X1 U1962 ( .C1(x1_ra_w[26]), .C2(n1098), .A(n1334), .B(n1335), .ZN(
        n1324) );
  AOI221_X1 U1963 ( .B1(x9_s1_w[27]), .B2(n1113), .C1(x8_s0_w[27]), .C2(n1114), 
        .A(n1321), .ZN(n1305) );
  AOI221_X1 U1964 ( .B1(x15_a5_w[27]), .B2(n1108), .C1(x14_a4_w[27]), .C2(
        n1109), .A(n1320), .ZN(n1306) );
  AOI211_X1 U1965 ( .C1(x1_ra_w[27]), .C2(n1098), .A(n1317), .B(n1318), .ZN(
        n1307) );
  AOI221_X1 U1966 ( .B1(x9_s1_w[28]), .B2(n1113), .C1(x8_s0_w[28]), .C2(n1114), 
        .A(n1304), .ZN(n1288) );
  AOI221_X1 U1967 ( .B1(x15_a5_w[28]), .B2(n1108), .C1(x14_a4_w[28]), .C2(
        n1109), .A(n1303), .ZN(n1289) );
  AOI211_X1 U1968 ( .C1(x1_ra_w[28]), .C2(n1098), .A(n1300), .B(n1301), .ZN(
        n1290) );
  AOI221_X1 U1969 ( .B1(x9_s1_w[29]), .B2(n1113), .C1(x8_s0_w[29]), .C2(n1114), 
        .A(n1287), .ZN(n1271) );
  AOI221_X1 U1970 ( .B1(x15_a5_w[29]), .B2(n1108), .C1(x14_a4_w[29]), .C2(
        n1109), .A(n1286), .ZN(n1272) );
  AOI211_X1 U1971 ( .C1(x1_ra_w[29]), .C2(n1098), .A(n1283), .B(n1284), .ZN(
        n1273) );
  AOI221_X1 U1972 ( .B1(x9_s1_w[30]), .B2(n1113), .C1(x8_s0_w[30]), .C2(n1114), 
        .A(n1253), .ZN(n1237) );
  AOI221_X1 U1973 ( .B1(x15_a5_w[30]), .B2(n1108), .C1(x14_a4_w[30]), .C2(
        n1109), .A(n1252), .ZN(n1238) );
  AOI211_X1 U1974 ( .C1(x1_ra_w[30]), .C2(n1098), .A(n1249), .B(n1250), .ZN(
        n1239) );
  AOI221_X1 U1975 ( .B1(x9_s1_w[31]), .B2(n1113), .C1(x8_s0_w[31]), .C2(n1114), 
        .A(n1236), .ZN(n1220) );
  AOI221_X1 U1976 ( .B1(x15_a5_w[31]), .B2(n1108), .C1(x14_a4_w[31]), .C2(
        n1109), .A(n1235), .ZN(n1221) );
  AOI211_X1 U1977 ( .C1(x1_ra_w[31]), .C2(n1098), .A(n1232), .B(n1233), .ZN(
        n1222) );
  AOI221_X1 U1978 ( .B1(n1703), .B2(x9_s1_w[0]), .C1(n1704), .C2(x8_s0_w[0]), 
        .A(n2248), .ZN(n2218) );
  AOI221_X1 U1979 ( .B1(n1698), .B2(x15_a5_w[0]), .C1(n1699), .C2(x14_a4_w[0]), 
        .A(n2247), .ZN(n2219) );
  AOI211_X1 U1980 ( .C1(n1688), .C2(x1_ra_w[0]), .A(n2240), .B(n2241), .ZN(
        n2220) );
  AOI221_X1 U1981 ( .B1(n1703), .B2(x9_s1_w[1]), .C1(n1704), .C2(x8_s0_w[1]), 
        .A(n2047), .ZN(n2031) );
  AOI221_X1 U1982 ( .B1(n1698), .B2(x15_a5_w[1]), .C1(n1699), .C2(x14_a4_w[1]), 
        .A(n2046), .ZN(n2032) );
  AOI211_X1 U1983 ( .C1(n1688), .C2(x1_ra_w[1]), .A(n2043), .B(n2044), .ZN(
        n2033) );
  AOI221_X1 U1984 ( .B1(n1703), .B2(x9_s1_w[2]), .C1(n1704), .C2(x8_s0_w[2]), 
        .A(n1860), .ZN(n1844) );
  AOI221_X1 U1985 ( .B1(n1698), .B2(x15_a5_w[2]), .C1(n1699), .C2(x14_a4_w[2]), 
        .A(n1859), .ZN(n1845) );
  AOI211_X1 U1986 ( .C1(n1688), .C2(x1_ra_w[2]), .A(n1856), .B(n1857), .ZN(
        n1846) );
  AOI221_X1 U1987 ( .B1(n1703), .B2(x9_s1_w[3]), .C1(n1704), .C2(x8_s0_w[3]), 
        .A(n1809), .ZN(n1793) );
  AOI221_X1 U1988 ( .B1(n1698), .B2(x15_a5_w[3]), .C1(n1699), .C2(x14_a4_w[3]), 
        .A(n1808), .ZN(n1794) );
  AOI211_X1 U1989 ( .C1(n1688), .C2(x1_ra_w[3]), .A(n1805), .B(n1806), .ZN(
        n1795) );
  AOI221_X1 U1990 ( .B1(n1703), .B2(x9_s1_w[4]), .C1(n1704), .C2(x8_s0_w[4]), 
        .A(n1792), .ZN(n1776) );
  AOI221_X1 U1991 ( .B1(n1698), .B2(x15_a5_w[4]), .C1(n1699), .C2(x14_a4_w[4]), 
        .A(n1791), .ZN(n1777) );
  AOI211_X1 U1992 ( .C1(n1688), .C2(x1_ra_w[4]), .A(n1788), .B(n1789), .ZN(
        n1778) );
  AOI221_X1 U1993 ( .B1(n1703), .B2(x9_s1_w[5]), .C1(n1704), .C2(x8_s0_w[5]), 
        .A(n1775), .ZN(n1759) );
  AOI221_X1 U1994 ( .B1(n1698), .B2(x15_a5_w[5]), .C1(n1699), .C2(x14_a4_w[5]), 
        .A(n1774), .ZN(n1760) );
  AOI211_X1 U1995 ( .C1(n1688), .C2(x1_ra_w[5]), .A(n1771), .B(n1772), .ZN(
        n1761) );
  AOI221_X1 U1996 ( .B1(n1703), .B2(x9_s1_w[6]), .C1(n1704), .C2(x8_s0_w[6]), 
        .A(n1758), .ZN(n1742) );
  AOI221_X1 U1997 ( .B1(n1698), .B2(x15_a5_w[6]), .C1(n1699), .C2(x14_a4_w[6]), 
        .A(n1757), .ZN(n1743) );
  AOI211_X1 U1998 ( .C1(n1688), .C2(x1_ra_w[6]), .A(n1754), .B(n1755), .ZN(
        n1744) );
  AOI221_X1 U1999 ( .B1(n1703), .B2(x9_s1_w[7]), .C1(n1704), .C2(x8_s0_w[7]), 
        .A(n1741), .ZN(n1725) );
  AOI221_X1 U2000 ( .B1(n1698), .B2(x15_a5_w[7]), .C1(n1699), .C2(x14_a4_w[7]), 
        .A(n1740), .ZN(n1726) );
  AOI211_X1 U2001 ( .C1(n1688), .C2(x1_ra_w[7]), .A(n1737), .B(n1738), .ZN(
        n1727) );
  AOI221_X1 U2002 ( .B1(n1703), .B2(x9_s1_w[8]), .C1(n1704), .C2(x8_s0_w[8]), 
        .A(n1724), .ZN(n1708) );
  AOI221_X1 U2003 ( .B1(n1698), .B2(x15_a5_w[8]), .C1(n1699), .C2(x14_a4_w[8]), 
        .A(n1723), .ZN(n1709) );
  AOI211_X1 U2004 ( .C1(n1688), .C2(x1_ra_w[8]), .A(n1720), .B(n1721), .ZN(
        n1710) );
  AOI221_X1 U2005 ( .B1(n1703), .B2(x9_s1_w[9]), .C1(n1704), .C2(x8_s0_w[9]), 
        .A(n1705), .ZN(n1660) );
  AOI221_X1 U2006 ( .B1(n1698), .B2(x15_a5_w[9]), .C1(n1699), .C2(x14_a4_w[9]), 
        .A(n1700), .ZN(n1661) );
  AOI211_X1 U2007 ( .C1(n1688), .C2(x1_ra_w[9]), .A(n1689), .B(n1690), .ZN(
        n1662) );
  AOI221_X1 U2008 ( .B1(n1703), .B2(x9_s1_w[10]), .C1(n1704), .C2(x8_s0_w[10]), 
        .A(n2217), .ZN(n2201) );
  AOI221_X1 U2009 ( .B1(n1698), .B2(x15_a5_w[10]), .C1(n1699), .C2(
        x14_a4_w[10]), .A(n2216), .ZN(n2202) );
  AOI211_X1 U2010 ( .C1(n1688), .C2(x1_ra_w[10]), .A(n2213), .B(n2214), .ZN(
        n2203) );
  AOI221_X1 U2011 ( .B1(n1703), .B2(x9_s1_w[11]), .C1(n1704), .C2(x8_s0_w[11]), 
        .A(n2200), .ZN(n2184) );
  AOI221_X1 U2012 ( .B1(n1698), .B2(x15_a5_w[11]), .C1(n1699), .C2(
        x14_a4_w[11]), .A(n2199), .ZN(n2185) );
  AOI211_X1 U2013 ( .C1(n1688), .C2(x1_ra_w[11]), .A(n2196), .B(n2197), .ZN(
        n2186) );
  AOI221_X1 U2014 ( .B1(n1703), .B2(x9_s1_w[12]), .C1(n1704), .C2(x8_s0_w[12]), 
        .A(n2183), .ZN(n2167) );
  AOI221_X1 U2015 ( .B1(n1698), .B2(x15_a5_w[12]), .C1(n1699), .C2(
        x14_a4_w[12]), .A(n2182), .ZN(n2168) );
  AOI211_X1 U2016 ( .C1(n1688), .C2(x1_ra_w[12]), .A(n2179), .B(n2180), .ZN(
        n2169) );
  AOI221_X1 U2017 ( .B1(n1703), .B2(x9_s1_w[13]), .C1(n1704), .C2(x8_s0_w[13]), 
        .A(n2166), .ZN(n2150) );
  AOI221_X1 U2018 ( .B1(n1698), .B2(x15_a5_w[13]), .C1(n1699), .C2(
        x14_a4_w[13]), .A(n2165), .ZN(n2151) );
  AOI211_X1 U2019 ( .C1(n1688), .C2(x1_ra_w[13]), .A(n2162), .B(n2163), .ZN(
        n2152) );
  AOI221_X1 U2020 ( .B1(n1703), .B2(x9_s1_w[14]), .C1(n1704), .C2(x8_s0_w[14]), 
        .A(n2149), .ZN(n2133) );
  AOI221_X1 U2021 ( .B1(n1698), .B2(x15_a5_w[14]), .C1(n1699), .C2(
        x14_a4_w[14]), .A(n2148), .ZN(n2134) );
  AOI211_X1 U2022 ( .C1(n1688), .C2(x1_ra_w[14]), .A(n2145), .B(n2146), .ZN(
        n2135) );
  AOI221_X1 U2023 ( .B1(n1703), .B2(x9_s1_w[15]), .C1(n1704), .C2(x8_s0_w[15]), 
        .A(n2132), .ZN(n2116) );
  AOI221_X1 U2024 ( .B1(n1698), .B2(x15_a5_w[15]), .C1(n1699), .C2(
        x14_a4_w[15]), .A(n2131), .ZN(n2117) );
  AOI211_X1 U2025 ( .C1(n1688), .C2(x1_ra_w[15]), .A(n2128), .B(n2129), .ZN(
        n2118) );
  AOI221_X1 U2026 ( .B1(n1703), .B2(x9_s1_w[16]), .C1(n1704), .C2(x8_s0_w[16]), 
        .A(n2115), .ZN(n2099) );
  AOI221_X1 U2027 ( .B1(n1698), .B2(x15_a5_w[16]), .C1(n1699), .C2(
        x14_a4_w[16]), .A(n2114), .ZN(n2100) );
  AOI211_X1 U2028 ( .C1(n1688), .C2(x1_ra_w[16]), .A(n2111), .B(n2112), .ZN(
        n2101) );
  AOI221_X1 U2029 ( .B1(n1703), .B2(x9_s1_w[17]), .C1(n1704), .C2(x8_s0_w[17]), 
        .A(n2098), .ZN(n2082) );
  AOI221_X1 U2030 ( .B1(n1698), .B2(x15_a5_w[17]), .C1(n1699), .C2(
        x14_a4_w[17]), .A(n2097), .ZN(n2083) );
  AOI211_X1 U2031 ( .C1(n1688), .C2(x1_ra_w[17]), .A(n2094), .B(n2095), .ZN(
        n2084) );
  AOI221_X1 U2032 ( .B1(n1703), .B2(x9_s1_w[18]), .C1(n1704), .C2(x8_s0_w[18]), 
        .A(n2081), .ZN(n2065) );
  AOI221_X1 U2033 ( .B1(n1698), .B2(x15_a5_w[18]), .C1(n1699), .C2(
        x14_a4_w[18]), .A(n2080), .ZN(n2066) );
  AOI211_X1 U2034 ( .C1(n1688), .C2(x1_ra_w[18]), .A(n2077), .B(n2078), .ZN(
        n2067) );
  AOI221_X1 U2035 ( .B1(n1703), .B2(x9_s1_w[19]), .C1(n1704), .C2(x8_s0_w[19]), 
        .A(n2064), .ZN(n2048) );
  AOI221_X1 U2036 ( .B1(n1698), .B2(x15_a5_w[19]), .C1(n1699), .C2(
        x14_a4_w[19]), .A(n2063), .ZN(n2049) );
  AOI211_X1 U2037 ( .C1(n1688), .C2(x1_ra_w[19]), .A(n2060), .B(n2061), .ZN(
        n2050) );
  AOI221_X1 U2038 ( .B1(n1703), .B2(x9_s1_w[20]), .C1(n1704), .C2(x8_s0_w[20]), 
        .A(n2030), .ZN(n2014) );
  AOI221_X1 U2039 ( .B1(n1698), .B2(x15_a5_w[20]), .C1(n1699), .C2(
        x14_a4_w[20]), .A(n2029), .ZN(n2015) );
  AOI211_X1 U2040 ( .C1(n1688), .C2(x1_ra_w[20]), .A(n2026), .B(n2027), .ZN(
        n2016) );
  AOI221_X1 U2041 ( .B1(n1703), .B2(x9_s1_w[21]), .C1(n1704), .C2(x8_s0_w[21]), 
        .A(n2013), .ZN(n1997) );
  AOI221_X1 U2042 ( .B1(n1698), .B2(x15_a5_w[21]), .C1(n1699), .C2(
        x14_a4_w[21]), .A(n2012), .ZN(n1998) );
  AOI211_X1 U2043 ( .C1(n1688), .C2(x1_ra_w[21]), .A(n2009), .B(n2010), .ZN(
        n1999) );
  AOI221_X1 U2044 ( .B1(n1703), .B2(x9_s1_w[22]), .C1(n1704), .C2(x8_s0_w[22]), 
        .A(n1996), .ZN(n1980) );
  AOI221_X1 U2045 ( .B1(n1698), .B2(x15_a5_w[22]), .C1(n1699), .C2(
        x14_a4_w[22]), .A(n1995), .ZN(n1981) );
  AOI211_X1 U2046 ( .C1(n1688), .C2(x1_ra_w[22]), .A(n1992), .B(n1993), .ZN(
        n1982) );
  AOI221_X1 U2047 ( .B1(n1703), .B2(x9_s1_w[23]), .C1(n1704), .C2(x8_s0_w[23]), 
        .A(n1979), .ZN(n1963) );
  AOI221_X1 U2048 ( .B1(n1698), .B2(x15_a5_w[23]), .C1(n1699), .C2(
        x14_a4_w[23]), .A(n1978), .ZN(n1964) );
  AOI211_X1 U2049 ( .C1(n1688), .C2(x1_ra_w[23]), .A(n1975), .B(n1976), .ZN(
        n1965) );
  AOI221_X1 U2050 ( .B1(n1703), .B2(x9_s1_w[24]), .C1(n1704), .C2(x8_s0_w[24]), 
        .A(n1962), .ZN(n1946) );
  AOI221_X1 U2051 ( .B1(n1698), .B2(x15_a5_w[24]), .C1(n1699), .C2(
        x14_a4_w[24]), .A(n1961), .ZN(n1947) );
  AOI211_X1 U2052 ( .C1(n1688), .C2(x1_ra_w[24]), .A(n1958), .B(n1959), .ZN(
        n1948) );
  AOI221_X1 U2053 ( .B1(n1703), .B2(x9_s1_w[25]), .C1(n1704), .C2(x8_s0_w[25]), 
        .A(n1945), .ZN(n1929) );
  AOI221_X1 U2054 ( .B1(n1698), .B2(x15_a5_w[25]), .C1(n1699), .C2(
        x14_a4_w[25]), .A(n1944), .ZN(n1930) );
  AOI211_X1 U2055 ( .C1(n1688), .C2(x1_ra_w[25]), .A(n1941), .B(n1942), .ZN(
        n1931) );
  AOI221_X1 U2056 ( .B1(n1703), .B2(x9_s1_w[26]), .C1(n1704), .C2(x8_s0_w[26]), 
        .A(n1928), .ZN(n1912) );
  AOI221_X1 U2057 ( .B1(n1698), .B2(x15_a5_w[26]), .C1(n1699), .C2(
        x14_a4_w[26]), .A(n1927), .ZN(n1913) );
  AOI211_X1 U2058 ( .C1(n1688), .C2(x1_ra_w[26]), .A(n1924), .B(n1925), .ZN(
        n1914) );
  AOI221_X1 U2059 ( .B1(n1703), .B2(x9_s1_w[27]), .C1(n1704), .C2(x8_s0_w[27]), 
        .A(n1911), .ZN(n1895) );
  AOI221_X1 U2060 ( .B1(n1698), .B2(x15_a5_w[27]), .C1(n1699), .C2(
        x14_a4_w[27]), .A(n1910), .ZN(n1896) );
  AOI211_X1 U2061 ( .C1(n1688), .C2(x1_ra_w[27]), .A(n1907), .B(n1908), .ZN(
        n1897) );
  AOI221_X1 U2062 ( .B1(n1703), .B2(x9_s1_w[28]), .C1(n1704), .C2(x8_s0_w[28]), 
        .A(n1894), .ZN(n1878) );
  AOI221_X1 U2063 ( .B1(n1698), .B2(x15_a5_w[28]), .C1(n1699), .C2(
        x14_a4_w[28]), .A(n1893), .ZN(n1879) );
  AOI211_X1 U2064 ( .C1(n1688), .C2(x1_ra_w[28]), .A(n1890), .B(n1891), .ZN(
        n1880) );
  AOI221_X1 U2065 ( .B1(n1703), .B2(x9_s1_w[29]), .C1(n1704), .C2(x8_s0_w[29]), 
        .A(n1877), .ZN(n1861) );
  AOI221_X1 U2066 ( .B1(n1698), .B2(x15_a5_w[29]), .C1(n1699), .C2(
        x14_a4_w[29]), .A(n1876), .ZN(n1862) );
  AOI211_X1 U2067 ( .C1(n1688), .C2(x1_ra_w[29]), .A(n1873), .B(n1874), .ZN(
        n1863) );
  AOI221_X1 U2068 ( .B1(n1703), .B2(x9_s1_w[30]), .C1(n1704), .C2(x8_s0_w[30]), 
        .A(n1843), .ZN(n1827) );
  AOI221_X1 U2069 ( .B1(n1698), .B2(x15_a5_w[30]), .C1(n1699), .C2(
        x14_a4_w[30]), .A(n1842), .ZN(n1828) );
  AOI211_X1 U2070 ( .C1(n1688), .C2(x1_ra_w[30]), .A(n1839), .B(n1840), .ZN(
        n1829) );
  AOI221_X1 U2071 ( .B1(n1703), .B2(x9_s1_w[31]), .C1(n1704), .C2(x8_s0_w[31]), 
        .A(n1826), .ZN(n1810) );
  AOI221_X1 U2072 ( .B1(n1698), .B2(x15_a5_w[31]), .C1(n1699), .C2(
        x14_a4_w[31]), .A(n1825), .ZN(n1811) );
  AOI211_X1 U2073 ( .C1(n1688), .C2(x1_ra_w[31]), .A(n1822), .B(n1823), .ZN(
        n1812) );
  AND2_X1 U2074 ( .A1(wa[4]), .A2(en_write), .ZN(n2360) );
  INV_X1 U2075 ( .A(wa[2]), .ZN(n3712) );
  INV_X1 U2076 ( .A(wa[0]), .ZN(n3714) );
  INV_X1 U2077 ( .A(wa[3]), .ZN(n3711) );
  INV_X1 U2078 ( .A(wa[1]), .ZN(n3713) );
  INV_X1 U2079 ( .A(n2289), .ZN(n3709) );
  AOI22_X1 U2080 ( .A1(wdata[0]), .A2(n581), .B1(n2290), .B2(x23_s7_w[0]), 
        .ZN(n2289) );
  INV_X1 U2081 ( .A(n2291), .ZN(n3693) );
  AOI22_X1 U2082 ( .A1(wdata[1]), .A2(n580), .B1(n2290), .B2(x23_s7_w[1]), 
        .ZN(n2291) );
  INV_X1 U2083 ( .A(n2292), .ZN(n3677) );
  AOI22_X1 U2084 ( .A1(wdata[2]), .A2(n581), .B1(n2290), .B2(x23_s7_w[2]), 
        .ZN(n2292) );
  INV_X1 U2085 ( .A(n2293), .ZN(n3661) );
  AOI22_X1 U2086 ( .A1(wdata[3]), .A2(n580), .B1(n2290), .B2(x23_s7_w[3]), 
        .ZN(n2293) );
  INV_X1 U2087 ( .A(n2294), .ZN(n3645) );
  AOI22_X1 U2088 ( .A1(wdata[4]), .A2(n581), .B1(n2290), .B2(x23_s7_w[4]), 
        .ZN(n2294) );
  INV_X1 U2089 ( .A(n2295), .ZN(n3629) );
  AOI22_X1 U2090 ( .A1(wdata[5]), .A2(n580), .B1(n2290), .B2(x23_s7_w[5]), 
        .ZN(n2295) );
  INV_X1 U2091 ( .A(n2296), .ZN(n3613) );
  AOI22_X1 U2092 ( .A1(wdata[6]), .A2(n581), .B1(n2290), .B2(x23_s7_w[6]), 
        .ZN(n2296) );
  INV_X1 U2093 ( .A(n2297), .ZN(n3597) );
  AOI22_X1 U2094 ( .A1(wdata[7]), .A2(n580), .B1(n2290), .B2(x23_s7_w[7]), 
        .ZN(n2297) );
  INV_X1 U2095 ( .A(n2298), .ZN(n3581) );
  AOI22_X1 U2096 ( .A1(wdata[8]), .A2(n581), .B1(n2290), .B2(x23_s7_w[8]), 
        .ZN(n2298) );
  INV_X1 U2097 ( .A(n2299), .ZN(n3565) );
  AOI22_X1 U2098 ( .A1(wdata[9]), .A2(n581), .B1(n2290), .B2(x23_s7_w[9]), 
        .ZN(n2299) );
  INV_X1 U2099 ( .A(n2300), .ZN(n3549) );
  AOI22_X1 U2100 ( .A1(wdata[10]), .A2(n581), .B1(n2290), .B2(x23_s7_w[10]), 
        .ZN(n2300) );
  INV_X1 U2101 ( .A(n2301), .ZN(n3533) );
  AOI22_X1 U2102 ( .A1(wdata[11]), .A2(n581), .B1(n2290), .B2(x23_s7_w[11]), 
        .ZN(n2301) );
  INV_X1 U2103 ( .A(n2302), .ZN(n3517) );
  AOI22_X1 U2104 ( .A1(wdata[12]), .A2(n581), .B1(n2290), .B2(x23_s7_w[12]), 
        .ZN(n2302) );
  INV_X1 U2105 ( .A(n2303), .ZN(n3501) );
  AOI22_X1 U2106 ( .A1(wdata[13]), .A2(n581), .B1(n2290), .B2(x23_s7_w[13]), 
        .ZN(n2303) );
  INV_X1 U2107 ( .A(n2304), .ZN(n3485) );
  AOI22_X1 U2108 ( .A1(wdata[14]), .A2(n581), .B1(n2290), .B2(x23_s7_w[14]), 
        .ZN(n2304) );
  INV_X1 U2109 ( .A(n2305), .ZN(n3469) );
  AOI22_X1 U2110 ( .A1(wdata[15]), .A2(n581), .B1(n2290), .B2(x23_s7_w[15]), 
        .ZN(n2305) );
  INV_X1 U2111 ( .A(n2306), .ZN(n3453) );
  AOI22_X1 U2112 ( .A1(wdata[16]), .A2(n581), .B1(n2290), .B2(x23_s7_w[16]), 
        .ZN(n2306) );
  INV_X1 U2113 ( .A(n2307), .ZN(n3437) );
  AOI22_X1 U2114 ( .A1(wdata[17]), .A2(n581), .B1(n2290), .B2(x23_s7_w[17]), 
        .ZN(n2307) );
  INV_X1 U2115 ( .A(n2308), .ZN(n3421) );
  AOI22_X1 U2116 ( .A1(wdata[18]), .A2(n581), .B1(n2290), .B2(x23_s7_w[18]), 
        .ZN(n2308) );
  INV_X1 U2117 ( .A(n2309), .ZN(n3405) );
  AOI22_X1 U2118 ( .A1(wdata[19]), .A2(n581), .B1(n2290), .B2(x23_s7_w[19]), 
        .ZN(n2309) );
  INV_X1 U2119 ( .A(n2310), .ZN(n3389) );
  AOI22_X1 U2120 ( .A1(wdata[20]), .A2(n580), .B1(n2290), .B2(x23_s7_w[20]), 
        .ZN(n2310) );
  INV_X1 U2121 ( .A(n2311), .ZN(n3373) );
  AOI22_X1 U2122 ( .A1(wdata[21]), .A2(n580), .B1(n2290), .B2(x23_s7_w[21]), 
        .ZN(n2311) );
  INV_X1 U2123 ( .A(n2312), .ZN(n3357) );
  AOI22_X1 U2124 ( .A1(wdata[22]), .A2(n580), .B1(n2290), .B2(x23_s7_w[22]), 
        .ZN(n2312) );
  INV_X1 U2125 ( .A(n2313), .ZN(n3341) );
  AOI22_X1 U2126 ( .A1(wdata[23]), .A2(n580), .B1(n2290), .B2(x23_s7_w[23]), 
        .ZN(n2313) );
  INV_X1 U2127 ( .A(n2314), .ZN(n3325) );
  AOI22_X1 U2128 ( .A1(wdata[24]), .A2(n580), .B1(n2290), .B2(x23_s7_w[24]), 
        .ZN(n2314) );
  INV_X1 U2129 ( .A(n2315), .ZN(n3309) );
  AOI22_X1 U2130 ( .A1(wdata[25]), .A2(n580), .B1(n2290), .B2(x23_s7_w[25]), 
        .ZN(n2315) );
  INV_X1 U2131 ( .A(n2316), .ZN(n3293) );
  AOI22_X1 U2132 ( .A1(wdata[26]), .A2(n580), .B1(n2290), .B2(x23_s7_w[26]), 
        .ZN(n2316) );
  INV_X1 U2133 ( .A(n2317), .ZN(n2357) );
  AOI22_X1 U2134 ( .A1(wdata[27]), .A2(n580), .B1(n2290), .B2(x23_s7_w[27]), 
        .ZN(n2317) );
  INV_X1 U2135 ( .A(n2318), .ZN(n1056) );
  AOI22_X1 U2136 ( .A1(wdata[28]), .A2(n580), .B1(n2290), .B2(x23_s7_w[28]), 
        .ZN(n2318) );
  INV_X1 U2137 ( .A(n2319), .ZN(n1040) );
  AOI22_X1 U2138 ( .A1(wdata[29]), .A2(n580), .B1(n2290), .B2(x23_s7_w[29]), 
        .ZN(n2319) );
  INV_X1 U2139 ( .A(n2320), .ZN(n1024) );
  AOI22_X1 U2140 ( .A1(wdata[30]), .A2(n580), .B1(n2290), .B2(x23_s7_w[30]), 
        .ZN(n2320) );
  INV_X1 U2141 ( .A(n2321), .ZN(n1008) );
  AOI22_X1 U2142 ( .A1(wdata[31]), .A2(n580), .B1(n2290), .B2(x23_s7_w[31]), 
        .ZN(n2321) );
  INV_X1 U2143 ( .A(n2324), .ZN(n3708) );
  AOI22_X1 U2144 ( .A1(wdata[0]), .A2(n444), .B1(n2325), .B2(x22_s6_w[0]), 
        .ZN(n2324) );
  INV_X1 U2145 ( .A(n2326), .ZN(n3692) );
  AOI22_X1 U2146 ( .A1(wdata[1]), .A2(n443), .B1(n2325), .B2(x22_s6_w[1]), 
        .ZN(n2326) );
  INV_X1 U2147 ( .A(n2327), .ZN(n3676) );
  AOI22_X1 U2148 ( .A1(wdata[2]), .A2(n444), .B1(n2325), .B2(x22_s6_w[2]), 
        .ZN(n2327) );
  INV_X1 U2149 ( .A(n2328), .ZN(n3660) );
  AOI22_X1 U2150 ( .A1(wdata[3]), .A2(n443), .B1(n2325), .B2(x22_s6_w[3]), 
        .ZN(n2328) );
  INV_X1 U2151 ( .A(n2329), .ZN(n3644) );
  AOI22_X1 U2152 ( .A1(wdata[4]), .A2(n444), .B1(n2325), .B2(x22_s6_w[4]), 
        .ZN(n2329) );
  INV_X1 U2153 ( .A(n2330), .ZN(n3628) );
  AOI22_X1 U2154 ( .A1(wdata[5]), .A2(n443), .B1(n2325), .B2(x22_s6_w[5]), 
        .ZN(n2330) );
  INV_X1 U2155 ( .A(n2331), .ZN(n3612) );
  AOI22_X1 U2156 ( .A1(wdata[6]), .A2(n444), .B1(n2325), .B2(x22_s6_w[6]), 
        .ZN(n2331) );
  INV_X1 U2157 ( .A(n2332), .ZN(n3596) );
  AOI22_X1 U2158 ( .A1(wdata[7]), .A2(n443), .B1(n2325), .B2(x22_s6_w[7]), 
        .ZN(n2332) );
  INV_X1 U2159 ( .A(n2333), .ZN(n3580) );
  AOI22_X1 U2160 ( .A1(wdata[8]), .A2(n444), .B1(n2325), .B2(x22_s6_w[8]), 
        .ZN(n2333) );
  INV_X1 U2161 ( .A(n2334), .ZN(n3564) );
  AOI22_X1 U2162 ( .A1(wdata[9]), .A2(n444), .B1(n2325), .B2(x22_s6_w[9]), 
        .ZN(n2334) );
  INV_X1 U2163 ( .A(n2335), .ZN(n3548) );
  AOI22_X1 U2164 ( .A1(wdata[10]), .A2(n444), .B1(n2325), .B2(x22_s6_w[10]), 
        .ZN(n2335) );
  INV_X1 U2165 ( .A(n2336), .ZN(n3532) );
  AOI22_X1 U2166 ( .A1(wdata[11]), .A2(n444), .B1(n2325), .B2(x22_s6_w[11]), 
        .ZN(n2336) );
  INV_X1 U2167 ( .A(n2337), .ZN(n3516) );
  AOI22_X1 U2168 ( .A1(wdata[12]), .A2(n444), .B1(n2325), .B2(x22_s6_w[12]), 
        .ZN(n2337) );
  INV_X1 U2169 ( .A(n2338), .ZN(n3500) );
  AOI22_X1 U2170 ( .A1(wdata[13]), .A2(n444), .B1(n2325), .B2(x22_s6_w[13]), 
        .ZN(n2338) );
  INV_X1 U2171 ( .A(n2339), .ZN(n3484) );
  AOI22_X1 U2172 ( .A1(wdata[14]), .A2(n444), .B1(n2325), .B2(x22_s6_w[14]), 
        .ZN(n2339) );
  INV_X1 U2173 ( .A(n2340), .ZN(n3468) );
  AOI22_X1 U2174 ( .A1(wdata[15]), .A2(n444), .B1(n2325), .B2(x22_s6_w[15]), 
        .ZN(n2340) );
  INV_X1 U2175 ( .A(n2341), .ZN(n3452) );
  AOI22_X1 U2176 ( .A1(wdata[16]), .A2(n444), .B1(n2325), .B2(x22_s6_w[16]), 
        .ZN(n2341) );
  INV_X1 U2177 ( .A(n2342), .ZN(n3436) );
  AOI22_X1 U2178 ( .A1(wdata[17]), .A2(n444), .B1(n2325), .B2(x22_s6_w[17]), 
        .ZN(n2342) );
  INV_X1 U2179 ( .A(n2343), .ZN(n3420) );
  AOI22_X1 U2180 ( .A1(wdata[18]), .A2(n444), .B1(n2325), .B2(x22_s6_w[18]), 
        .ZN(n2343) );
  INV_X1 U2181 ( .A(n2344), .ZN(n3404) );
  AOI22_X1 U2182 ( .A1(wdata[19]), .A2(n444), .B1(n2325), .B2(x22_s6_w[19]), 
        .ZN(n2344) );
  INV_X1 U2183 ( .A(n2345), .ZN(n3388) );
  AOI22_X1 U2184 ( .A1(wdata[20]), .A2(n443), .B1(n2325), .B2(x22_s6_w[20]), 
        .ZN(n2345) );
  INV_X1 U2185 ( .A(n2346), .ZN(n3372) );
  AOI22_X1 U2186 ( .A1(wdata[21]), .A2(n443), .B1(n2325), .B2(x22_s6_w[21]), 
        .ZN(n2346) );
  INV_X1 U2187 ( .A(n2347), .ZN(n3356) );
  AOI22_X1 U2188 ( .A1(wdata[22]), .A2(n443), .B1(n2325), .B2(x22_s6_w[22]), 
        .ZN(n2347) );
  INV_X1 U2189 ( .A(n2348), .ZN(n3340) );
  AOI22_X1 U2190 ( .A1(wdata[23]), .A2(n443), .B1(n2325), .B2(x22_s6_w[23]), 
        .ZN(n2348) );
  INV_X1 U2191 ( .A(n2349), .ZN(n3324) );
  AOI22_X1 U2192 ( .A1(wdata[24]), .A2(n443), .B1(n2325), .B2(x22_s6_w[24]), 
        .ZN(n2349) );
  INV_X1 U2193 ( .A(n2350), .ZN(n3308) );
  AOI22_X1 U2194 ( .A1(wdata[25]), .A2(n443), .B1(n2325), .B2(x22_s6_w[25]), 
        .ZN(n2350) );
  INV_X1 U2195 ( .A(n2351), .ZN(n3292) );
  AOI22_X1 U2196 ( .A1(wdata[26]), .A2(n443), .B1(n2325), .B2(x22_s6_w[26]), 
        .ZN(n2351) );
  INV_X1 U2197 ( .A(n2352), .ZN(n2287) );
  AOI22_X1 U2198 ( .A1(wdata[27]), .A2(n443), .B1(n2325), .B2(x22_s6_w[27]), 
        .ZN(n2352) );
  INV_X1 U2199 ( .A(n2353), .ZN(n1055) );
  AOI22_X1 U2200 ( .A1(wdata[28]), .A2(n443), .B1(n2325), .B2(x22_s6_w[28]), 
        .ZN(n2353) );
  INV_X1 U2201 ( .A(n2354), .ZN(n1039) );
  AOI22_X1 U2202 ( .A1(wdata[29]), .A2(n443), .B1(n2325), .B2(x22_s6_w[29]), 
        .ZN(n2354) );
  INV_X1 U2203 ( .A(n2355), .ZN(n1023) );
  AOI22_X1 U2204 ( .A1(wdata[30]), .A2(n443), .B1(n2325), .B2(x22_s6_w[30]), 
        .ZN(n2355) );
  INV_X1 U2205 ( .A(n2356), .ZN(n1007) );
  AOI22_X1 U2206 ( .A1(wdata[31]), .A2(n443), .B1(n2325), .B2(x22_s6_w[31]), 
        .ZN(n2356) );
  INV_X1 U2207 ( .A(n2364), .ZN(n3707) );
  AOI22_X1 U2208 ( .A1(wdata[0]), .A2(n399), .B1(n2365), .B2(x17_a7_w[0]), 
        .ZN(n2364) );
  INV_X1 U2209 ( .A(n2366), .ZN(n3691) );
  AOI22_X1 U2210 ( .A1(wdata[1]), .A2(n398), .B1(n2365), .B2(x17_a7_w[1]), 
        .ZN(n2366) );
  INV_X1 U2211 ( .A(n2367), .ZN(n3675) );
  AOI22_X1 U2212 ( .A1(wdata[2]), .A2(n399), .B1(n2365), .B2(x17_a7_w[2]), 
        .ZN(n2367) );
  INV_X1 U2213 ( .A(n2368), .ZN(n3659) );
  AOI22_X1 U2214 ( .A1(wdata[3]), .A2(n398), .B1(n2365), .B2(x17_a7_w[3]), 
        .ZN(n2368) );
  INV_X1 U2215 ( .A(n2369), .ZN(n3643) );
  AOI22_X1 U2216 ( .A1(wdata[4]), .A2(n399), .B1(n2365), .B2(x17_a7_w[4]), 
        .ZN(n2369) );
  INV_X1 U2217 ( .A(n2370), .ZN(n3627) );
  AOI22_X1 U2218 ( .A1(wdata[5]), .A2(n398), .B1(n2365), .B2(x17_a7_w[5]), 
        .ZN(n2370) );
  INV_X1 U2219 ( .A(n2371), .ZN(n3611) );
  AOI22_X1 U2220 ( .A1(wdata[6]), .A2(n399), .B1(n2365), .B2(x17_a7_w[6]), 
        .ZN(n2371) );
  INV_X1 U2221 ( .A(n2372), .ZN(n3595) );
  AOI22_X1 U2222 ( .A1(wdata[7]), .A2(n398), .B1(n2365), .B2(x17_a7_w[7]), 
        .ZN(n2372) );
  INV_X1 U2223 ( .A(n2373), .ZN(n3579) );
  AOI22_X1 U2224 ( .A1(wdata[8]), .A2(n399), .B1(n2365), .B2(x17_a7_w[8]), 
        .ZN(n2373) );
  INV_X1 U2225 ( .A(n2374), .ZN(n3563) );
  AOI22_X1 U2226 ( .A1(wdata[9]), .A2(n399), .B1(n2365), .B2(x17_a7_w[9]), 
        .ZN(n2374) );
  INV_X1 U2227 ( .A(n2375), .ZN(n3547) );
  AOI22_X1 U2228 ( .A1(wdata[10]), .A2(n399), .B1(n2365), .B2(x17_a7_w[10]), 
        .ZN(n2375) );
  INV_X1 U2229 ( .A(n2376), .ZN(n3531) );
  AOI22_X1 U2230 ( .A1(wdata[11]), .A2(n399), .B1(n2365), .B2(x17_a7_w[11]), 
        .ZN(n2376) );
  INV_X1 U2231 ( .A(n2377), .ZN(n3515) );
  AOI22_X1 U2232 ( .A1(wdata[12]), .A2(n399), .B1(n2365), .B2(x17_a7_w[12]), 
        .ZN(n2377) );
  INV_X1 U2233 ( .A(n2378), .ZN(n3499) );
  AOI22_X1 U2234 ( .A1(wdata[13]), .A2(n399), .B1(n2365), .B2(x17_a7_w[13]), 
        .ZN(n2378) );
  INV_X1 U2235 ( .A(n2379), .ZN(n3483) );
  AOI22_X1 U2236 ( .A1(wdata[14]), .A2(n399), .B1(n2365), .B2(x17_a7_w[14]), 
        .ZN(n2379) );
  INV_X1 U2237 ( .A(n2380), .ZN(n3467) );
  AOI22_X1 U2238 ( .A1(wdata[15]), .A2(n399), .B1(n2365), .B2(x17_a7_w[15]), 
        .ZN(n2380) );
  INV_X1 U2239 ( .A(n2381), .ZN(n3451) );
  AOI22_X1 U2240 ( .A1(wdata[16]), .A2(n399), .B1(n2365), .B2(x17_a7_w[16]), 
        .ZN(n2381) );
  INV_X1 U2241 ( .A(n2382), .ZN(n3435) );
  AOI22_X1 U2242 ( .A1(wdata[17]), .A2(n399), .B1(n2365), .B2(x17_a7_w[17]), 
        .ZN(n2382) );
  INV_X1 U2243 ( .A(n2383), .ZN(n3419) );
  AOI22_X1 U2244 ( .A1(wdata[18]), .A2(n399), .B1(n2365), .B2(x17_a7_w[18]), 
        .ZN(n2383) );
  INV_X1 U2245 ( .A(n2384), .ZN(n3403) );
  AOI22_X1 U2246 ( .A1(wdata[19]), .A2(n399), .B1(n2365), .B2(x17_a7_w[19]), 
        .ZN(n2384) );
  INV_X1 U2247 ( .A(n2385), .ZN(n3387) );
  AOI22_X1 U2248 ( .A1(wdata[20]), .A2(n398), .B1(n2365), .B2(x17_a7_w[20]), 
        .ZN(n2385) );
  INV_X1 U2249 ( .A(n2386), .ZN(n3371) );
  AOI22_X1 U2250 ( .A1(wdata[21]), .A2(n398), .B1(n2365), .B2(x17_a7_w[21]), 
        .ZN(n2386) );
  INV_X1 U2251 ( .A(n2387), .ZN(n3355) );
  AOI22_X1 U2252 ( .A1(wdata[22]), .A2(n398), .B1(n2365), .B2(x17_a7_w[22]), 
        .ZN(n2387) );
  INV_X1 U2253 ( .A(n2388), .ZN(n3339) );
  AOI22_X1 U2254 ( .A1(wdata[23]), .A2(n398), .B1(n2365), .B2(x17_a7_w[23]), 
        .ZN(n2388) );
  INV_X1 U2255 ( .A(n2389), .ZN(n3323) );
  AOI22_X1 U2256 ( .A1(wdata[24]), .A2(n398), .B1(n2365), .B2(x17_a7_w[24]), 
        .ZN(n2389) );
  INV_X1 U2257 ( .A(n2390), .ZN(n3307) );
  AOI22_X1 U2258 ( .A1(wdata[25]), .A2(n398), .B1(n2365), .B2(x17_a7_w[25]), 
        .ZN(n2390) );
  INV_X1 U2259 ( .A(n2391), .ZN(n3291) );
  AOI22_X1 U2260 ( .A1(wdata[26]), .A2(n398), .B1(n2365), .B2(x17_a7_w[26]), 
        .ZN(n2391) );
  INV_X1 U2261 ( .A(n2392), .ZN(n2285) );
  AOI22_X1 U2262 ( .A1(wdata[27]), .A2(n398), .B1(n2365), .B2(x17_a7_w[27]), 
        .ZN(n2392) );
  INV_X1 U2263 ( .A(n2393), .ZN(n1054) );
  AOI22_X1 U2264 ( .A1(wdata[28]), .A2(n398), .B1(n2365), .B2(x17_a7_w[28]), 
        .ZN(n2393) );
  INV_X1 U2265 ( .A(n2394), .ZN(n1038) );
  AOI22_X1 U2266 ( .A1(wdata[29]), .A2(n398), .B1(n2365), .B2(x17_a7_w[29]), 
        .ZN(n2394) );
  INV_X1 U2267 ( .A(n2395), .ZN(n1022) );
  AOI22_X1 U2268 ( .A1(wdata[30]), .A2(n398), .B1(n2365), .B2(x17_a7_w[30]), 
        .ZN(n2395) );
  INV_X1 U2269 ( .A(n2396), .ZN(n1006) );
  AOI22_X1 U2270 ( .A1(wdata[31]), .A2(n398), .B1(n2365), .B2(x17_a7_w[31]), 
        .ZN(n2396) );
  INV_X1 U2271 ( .A(n2397), .ZN(n3706) );
  AOI22_X1 U2272 ( .A1(wdata[0]), .A2(n390), .B1(n2398), .B2(x16_a6_w[0]), 
        .ZN(n2397) );
  INV_X1 U2273 ( .A(n2399), .ZN(n3690) );
  AOI22_X1 U2274 ( .A1(wdata[1]), .A2(n389), .B1(n2398), .B2(x16_a6_w[1]), 
        .ZN(n2399) );
  INV_X1 U2275 ( .A(n2400), .ZN(n3674) );
  AOI22_X1 U2276 ( .A1(wdata[2]), .A2(n390), .B1(n2398), .B2(x16_a6_w[2]), 
        .ZN(n2400) );
  INV_X1 U2277 ( .A(n2401), .ZN(n3658) );
  AOI22_X1 U2278 ( .A1(wdata[3]), .A2(n389), .B1(n2398), .B2(x16_a6_w[3]), 
        .ZN(n2401) );
  INV_X1 U2279 ( .A(n2402), .ZN(n3642) );
  AOI22_X1 U2280 ( .A1(wdata[4]), .A2(n390), .B1(n2398), .B2(x16_a6_w[4]), 
        .ZN(n2402) );
  INV_X1 U2281 ( .A(n2403), .ZN(n3626) );
  AOI22_X1 U2282 ( .A1(wdata[5]), .A2(n389), .B1(n2398), .B2(x16_a6_w[5]), 
        .ZN(n2403) );
  INV_X1 U2283 ( .A(n2404), .ZN(n3610) );
  AOI22_X1 U2284 ( .A1(wdata[6]), .A2(n390), .B1(n2398), .B2(x16_a6_w[6]), 
        .ZN(n2404) );
  INV_X1 U2285 ( .A(n2405), .ZN(n3594) );
  AOI22_X1 U2286 ( .A1(wdata[7]), .A2(n389), .B1(n2398), .B2(x16_a6_w[7]), 
        .ZN(n2405) );
  INV_X1 U2287 ( .A(n2431), .ZN(n3705) );
  AOI22_X1 U2288 ( .A1(wdata[0]), .A2(n381), .B1(n2432), .B2(x15_a5_w[0]), 
        .ZN(n2431) );
  INV_X1 U2289 ( .A(n2433), .ZN(n3689) );
  AOI22_X1 U2290 ( .A1(wdata[1]), .A2(n380), .B1(n2432), .B2(x15_a5_w[1]), 
        .ZN(n2433) );
  INV_X1 U2291 ( .A(n2434), .ZN(n3673) );
  AOI22_X1 U2292 ( .A1(wdata[2]), .A2(n381), .B1(n2432), .B2(x15_a5_w[2]), 
        .ZN(n2434) );
  INV_X1 U2293 ( .A(n2435), .ZN(n3657) );
  AOI22_X1 U2294 ( .A1(wdata[3]), .A2(n380), .B1(n2432), .B2(x15_a5_w[3]), 
        .ZN(n2435) );
  INV_X1 U2295 ( .A(n2436), .ZN(n3641) );
  AOI22_X1 U2296 ( .A1(wdata[4]), .A2(n381), .B1(n2432), .B2(x15_a5_w[4]), 
        .ZN(n2436) );
  INV_X1 U2297 ( .A(n2437), .ZN(n3625) );
  AOI22_X1 U2298 ( .A1(wdata[5]), .A2(n380), .B1(n2432), .B2(x15_a5_w[5]), 
        .ZN(n2437) );
  INV_X1 U2299 ( .A(n2438), .ZN(n3609) );
  AOI22_X1 U2300 ( .A1(wdata[6]), .A2(n381), .B1(n2432), .B2(x15_a5_w[6]), 
        .ZN(n2438) );
  INV_X1 U2301 ( .A(n2439), .ZN(n3593) );
  AOI22_X1 U2302 ( .A1(wdata[7]), .A2(n380), .B1(n2432), .B2(x15_a5_w[7]), 
        .ZN(n2439) );
  INV_X1 U2303 ( .A(n2440), .ZN(n3577) );
  AOI22_X1 U2304 ( .A1(wdata[8]), .A2(n381), .B1(n2432), .B2(x15_a5_w[8]), 
        .ZN(n2440) );
  INV_X1 U2305 ( .A(n2441), .ZN(n3561) );
  AOI22_X1 U2306 ( .A1(wdata[9]), .A2(n381), .B1(n2432), .B2(x15_a5_w[9]), 
        .ZN(n2441) );
  INV_X1 U2307 ( .A(n2442), .ZN(n3545) );
  AOI22_X1 U2308 ( .A1(wdata[10]), .A2(n381), .B1(n2432), .B2(x15_a5_w[10]), 
        .ZN(n2442) );
  INV_X1 U2309 ( .A(n2443), .ZN(n3529) );
  AOI22_X1 U2310 ( .A1(wdata[11]), .A2(n381), .B1(n2432), .B2(x15_a5_w[11]), 
        .ZN(n2443) );
  INV_X1 U2311 ( .A(n2444), .ZN(n3513) );
  AOI22_X1 U2312 ( .A1(wdata[12]), .A2(n381), .B1(n2432), .B2(x15_a5_w[12]), 
        .ZN(n2444) );
  INV_X1 U2313 ( .A(n2445), .ZN(n3497) );
  AOI22_X1 U2314 ( .A1(wdata[13]), .A2(n381), .B1(n2432), .B2(x15_a5_w[13]), 
        .ZN(n2445) );
  INV_X1 U2315 ( .A(n2446), .ZN(n3481) );
  AOI22_X1 U2316 ( .A1(wdata[14]), .A2(n381), .B1(n2432), .B2(x15_a5_w[14]), 
        .ZN(n2446) );
  INV_X1 U2317 ( .A(n2447), .ZN(n3465) );
  AOI22_X1 U2318 ( .A1(wdata[15]), .A2(n381), .B1(n2432), .B2(x15_a5_w[15]), 
        .ZN(n2447) );
  INV_X1 U2319 ( .A(n2448), .ZN(n3449) );
  AOI22_X1 U2320 ( .A1(wdata[16]), .A2(n381), .B1(n2432), .B2(x15_a5_w[16]), 
        .ZN(n2448) );
  INV_X1 U2321 ( .A(n2449), .ZN(n3433) );
  AOI22_X1 U2322 ( .A1(wdata[17]), .A2(n381), .B1(n2432), .B2(x15_a5_w[17]), 
        .ZN(n2449) );
  INV_X1 U2323 ( .A(n2450), .ZN(n3417) );
  AOI22_X1 U2324 ( .A1(wdata[18]), .A2(n381), .B1(n2432), .B2(x15_a5_w[18]), 
        .ZN(n2450) );
  INV_X1 U2325 ( .A(n2451), .ZN(n3401) );
  AOI22_X1 U2326 ( .A1(wdata[19]), .A2(n381), .B1(n2432), .B2(x15_a5_w[19]), 
        .ZN(n2451) );
  INV_X1 U2327 ( .A(n2452), .ZN(n3385) );
  AOI22_X1 U2328 ( .A1(wdata[20]), .A2(n380), .B1(n2432), .B2(x15_a5_w[20]), 
        .ZN(n2452) );
  INV_X1 U2329 ( .A(n2453), .ZN(n3369) );
  AOI22_X1 U2330 ( .A1(wdata[21]), .A2(n380), .B1(n2432), .B2(x15_a5_w[21]), 
        .ZN(n2453) );
  INV_X1 U2331 ( .A(n2454), .ZN(n3353) );
  AOI22_X1 U2332 ( .A1(wdata[22]), .A2(n380), .B1(n2432), .B2(x15_a5_w[22]), 
        .ZN(n2454) );
  INV_X1 U2333 ( .A(n2455), .ZN(n3337) );
  AOI22_X1 U2334 ( .A1(wdata[23]), .A2(n380), .B1(n2432), .B2(x15_a5_w[23]), 
        .ZN(n2455) );
  INV_X1 U2335 ( .A(n2456), .ZN(n3321) );
  AOI22_X1 U2336 ( .A1(wdata[24]), .A2(n380), .B1(n2432), .B2(x15_a5_w[24]), 
        .ZN(n2456) );
  INV_X1 U2337 ( .A(n2457), .ZN(n3305) );
  AOI22_X1 U2338 ( .A1(wdata[25]), .A2(n380), .B1(n2432), .B2(x15_a5_w[25]), 
        .ZN(n2457) );
  INV_X1 U2339 ( .A(n2458), .ZN(n2777) );
  AOI22_X1 U2340 ( .A1(wdata[26]), .A2(n380), .B1(n2432), .B2(x15_a5_w[26]), 
        .ZN(n2458) );
  INV_X1 U2341 ( .A(n2459), .ZN(n1068) );
  AOI22_X1 U2342 ( .A1(wdata[27]), .A2(n380), .B1(n2432), .B2(x15_a5_w[27]), 
        .ZN(n2459) );
  INV_X1 U2343 ( .A(n2460), .ZN(n1052) );
  AOI22_X1 U2344 ( .A1(wdata[28]), .A2(n380), .B1(n2432), .B2(x15_a5_w[28]), 
        .ZN(n2460) );
  INV_X1 U2345 ( .A(n2461), .ZN(n1036) );
  AOI22_X1 U2346 ( .A1(wdata[29]), .A2(n380), .B1(n2432), .B2(x15_a5_w[29]), 
        .ZN(n2461) );
  INV_X1 U2347 ( .A(n2462), .ZN(n1020) );
  AOI22_X1 U2348 ( .A1(wdata[30]), .A2(n380), .B1(n2432), .B2(x15_a5_w[30]), 
        .ZN(n2462) );
  INV_X1 U2349 ( .A(n2463), .ZN(n1004) );
  AOI22_X1 U2350 ( .A1(wdata[31]), .A2(n380), .B1(n2432), .B2(x15_a5_w[31]), 
        .ZN(n2463) );
  INV_X1 U2351 ( .A(n2465), .ZN(n3704) );
  AOI22_X1 U2352 ( .A1(wdata[0]), .A2(n372), .B1(n2466), .B2(x14_a4_w[0]), 
        .ZN(n2465) );
  INV_X1 U2353 ( .A(n2467), .ZN(n3688) );
  AOI22_X1 U2354 ( .A1(wdata[1]), .A2(n371), .B1(n2466), .B2(x14_a4_w[1]), 
        .ZN(n2467) );
  INV_X1 U2355 ( .A(n2468), .ZN(n3672) );
  AOI22_X1 U2356 ( .A1(wdata[2]), .A2(n372), .B1(n2466), .B2(x14_a4_w[2]), 
        .ZN(n2468) );
  INV_X1 U2357 ( .A(n2469), .ZN(n3656) );
  AOI22_X1 U2358 ( .A1(wdata[3]), .A2(n371), .B1(n2466), .B2(x14_a4_w[3]), 
        .ZN(n2469) );
  INV_X1 U2359 ( .A(n2470), .ZN(n3640) );
  AOI22_X1 U2360 ( .A1(wdata[4]), .A2(n372), .B1(n2466), .B2(x14_a4_w[4]), 
        .ZN(n2470) );
  INV_X1 U2361 ( .A(n2471), .ZN(n3624) );
  AOI22_X1 U2362 ( .A1(wdata[5]), .A2(n371), .B1(n2466), .B2(x14_a4_w[5]), 
        .ZN(n2471) );
  INV_X1 U2363 ( .A(n2472), .ZN(n3608) );
  AOI22_X1 U2364 ( .A1(wdata[6]), .A2(n372), .B1(n2466), .B2(x14_a4_w[6]), 
        .ZN(n2472) );
  INV_X1 U2365 ( .A(n2473), .ZN(n3592) );
  AOI22_X1 U2366 ( .A1(wdata[7]), .A2(n371), .B1(n2466), .B2(x14_a4_w[7]), 
        .ZN(n2473) );
  INV_X1 U2367 ( .A(n2474), .ZN(n3576) );
  AOI22_X1 U2368 ( .A1(wdata[8]), .A2(n372), .B1(n2466), .B2(x14_a4_w[8]), 
        .ZN(n2474) );
  INV_X1 U2369 ( .A(n2475), .ZN(n3560) );
  AOI22_X1 U2370 ( .A1(wdata[9]), .A2(n372), .B1(n2466), .B2(x14_a4_w[9]), 
        .ZN(n2475) );
  INV_X1 U2371 ( .A(n2476), .ZN(n3544) );
  AOI22_X1 U2372 ( .A1(wdata[10]), .A2(n372), .B1(n2466), .B2(x14_a4_w[10]), 
        .ZN(n2476) );
  INV_X1 U2373 ( .A(n2477), .ZN(n3528) );
  AOI22_X1 U2374 ( .A1(wdata[11]), .A2(n372), .B1(n2466), .B2(x14_a4_w[11]), 
        .ZN(n2477) );
  INV_X1 U2375 ( .A(n2478), .ZN(n3512) );
  AOI22_X1 U2376 ( .A1(wdata[12]), .A2(n372), .B1(n2466), .B2(x14_a4_w[12]), 
        .ZN(n2478) );
  INV_X1 U2377 ( .A(n2479), .ZN(n3496) );
  AOI22_X1 U2378 ( .A1(wdata[13]), .A2(n372), .B1(n2466), .B2(x14_a4_w[13]), 
        .ZN(n2479) );
  INV_X1 U2379 ( .A(n2480), .ZN(n3480) );
  AOI22_X1 U2380 ( .A1(wdata[14]), .A2(n372), .B1(n2466), .B2(x14_a4_w[14]), 
        .ZN(n2480) );
  INV_X1 U2381 ( .A(n2481), .ZN(n3464) );
  AOI22_X1 U2382 ( .A1(wdata[15]), .A2(n372), .B1(n2466), .B2(x14_a4_w[15]), 
        .ZN(n2481) );
  INV_X1 U2383 ( .A(n2482), .ZN(n3448) );
  AOI22_X1 U2384 ( .A1(wdata[16]), .A2(n372), .B1(n2466), .B2(x14_a4_w[16]), 
        .ZN(n2482) );
  INV_X1 U2385 ( .A(n2483), .ZN(n3432) );
  AOI22_X1 U2386 ( .A1(wdata[17]), .A2(n372), .B1(n2466), .B2(x14_a4_w[17]), 
        .ZN(n2483) );
  INV_X1 U2387 ( .A(n2484), .ZN(n3416) );
  AOI22_X1 U2388 ( .A1(wdata[18]), .A2(n372), .B1(n2466), .B2(x14_a4_w[18]), 
        .ZN(n2484) );
  INV_X1 U2389 ( .A(n2485), .ZN(n3400) );
  AOI22_X1 U2390 ( .A1(wdata[19]), .A2(n372), .B1(n2466), .B2(x14_a4_w[19]), 
        .ZN(n2485) );
  INV_X1 U2391 ( .A(n2486), .ZN(n3384) );
  AOI22_X1 U2392 ( .A1(wdata[20]), .A2(n371), .B1(n2466), .B2(x14_a4_w[20]), 
        .ZN(n2486) );
  INV_X1 U2393 ( .A(n2487), .ZN(n3368) );
  AOI22_X1 U2394 ( .A1(wdata[21]), .A2(n371), .B1(n2466), .B2(x14_a4_w[21]), 
        .ZN(n2487) );
  INV_X1 U2395 ( .A(n2488), .ZN(n3352) );
  AOI22_X1 U2396 ( .A1(wdata[22]), .A2(n371), .B1(n2466), .B2(x14_a4_w[22]), 
        .ZN(n2488) );
  INV_X1 U2397 ( .A(n2489), .ZN(n3336) );
  AOI22_X1 U2398 ( .A1(wdata[23]), .A2(n371), .B1(n2466), .B2(x14_a4_w[23]), 
        .ZN(n2489) );
  INV_X1 U2399 ( .A(n2490), .ZN(n3320) );
  AOI22_X1 U2400 ( .A1(wdata[24]), .A2(n371), .B1(n2466), .B2(x14_a4_w[24]), 
        .ZN(n2490) );
  INV_X1 U2401 ( .A(n2491), .ZN(n3304) );
  AOI22_X1 U2402 ( .A1(wdata[25]), .A2(n371), .B1(n2466), .B2(x14_a4_w[25]), 
        .ZN(n2491) );
  INV_X1 U2403 ( .A(n2492), .ZN(n2643) );
  AOI22_X1 U2404 ( .A1(wdata[26]), .A2(n371), .B1(n2466), .B2(x14_a4_w[26]), 
        .ZN(n2492) );
  INV_X1 U2405 ( .A(n2493), .ZN(n1067) );
  AOI22_X1 U2406 ( .A1(wdata[27]), .A2(n371), .B1(n2466), .B2(x14_a4_w[27]), 
        .ZN(n2493) );
  INV_X1 U2407 ( .A(n2494), .ZN(n1051) );
  AOI22_X1 U2408 ( .A1(wdata[28]), .A2(n371), .B1(n2466), .B2(x14_a4_w[28]), 
        .ZN(n2494) );
  INV_X1 U2409 ( .A(n2495), .ZN(n1035) );
  AOI22_X1 U2410 ( .A1(wdata[29]), .A2(n371), .B1(n2466), .B2(x14_a4_w[29]), 
        .ZN(n2495) );
  INV_X1 U2411 ( .A(n2496), .ZN(n1019) );
  AOI22_X1 U2412 ( .A1(wdata[30]), .A2(n371), .B1(n2466), .B2(x14_a4_w[30]), 
        .ZN(n2496) );
  INV_X1 U2413 ( .A(n2497), .ZN(n1003) );
  AOI22_X1 U2414 ( .A1(wdata[31]), .A2(n371), .B1(n2466), .B2(x14_a4_w[31]), 
        .ZN(n2497) );
  INV_X1 U2415 ( .A(n2505), .ZN(n3703) );
  AOI22_X1 U2416 ( .A1(wdata[0]), .A2(n327), .B1(n2506), .B2(x9_s1_w[0]), .ZN(
        n2505) );
  INV_X1 U2417 ( .A(n2507), .ZN(n3687) );
  AOI22_X1 U2418 ( .A1(wdata[1]), .A2(n326), .B1(n2506), .B2(x9_s1_w[1]), .ZN(
        n2507) );
  INV_X1 U2419 ( .A(n2508), .ZN(n3671) );
  AOI22_X1 U2420 ( .A1(wdata[2]), .A2(n327), .B1(n2506), .B2(x9_s1_w[2]), .ZN(
        n2508) );
  INV_X1 U2421 ( .A(n2509), .ZN(n3655) );
  AOI22_X1 U2422 ( .A1(wdata[3]), .A2(n326), .B1(n2506), .B2(x9_s1_w[3]), .ZN(
        n2509) );
  INV_X1 U2423 ( .A(n2510), .ZN(n3639) );
  AOI22_X1 U2424 ( .A1(wdata[4]), .A2(n327), .B1(n2506), .B2(x9_s1_w[4]), .ZN(
        n2510) );
  INV_X1 U2425 ( .A(n2511), .ZN(n3623) );
  AOI22_X1 U2426 ( .A1(wdata[5]), .A2(n326), .B1(n2506), .B2(x9_s1_w[5]), .ZN(
        n2511) );
  INV_X1 U2427 ( .A(n2512), .ZN(n3607) );
  AOI22_X1 U2428 ( .A1(wdata[6]), .A2(n327), .B1(n2506), .B2(x9_s1_w[6]), .ZN(
        n2512) );
  INV_X1 U2429 ( .A(n2513), .ZN(n3591) );
  AOI22_X1 U2430 ( .A1(wdata[7]), .A2(n326), .B1(n2506), .B2(x9_s1_w[7]), .ZN(
        n2513) );
  INV_X1 U2431 ( .A(n2514), .ZN(n3575) );
  AOI22_X1 U2432 ( .A1(wdata[8]), .A2(n327), .B1(n2506), .B2(x9_s1_w[8]), .ZN(
        n2514) );
  INV_X1 U2433 ( .A(n2515), .ZN(n3559) );
  AOI22_X1 U2434 ( .A1(wdata[9]), .A2(n327), .B1(n2506), .B2(x9_s1_w[9]), .ZN(
        n2515) );
  INV_X1 U2435 ( .A(n2516), .ZN(n3543) );
  AOI22_X1 U2436 ( .A1(wdata[10]), .A2(n327), .B1(n2506), .B2(x9_s1_w[10]), 
        .ZN(n2516) );
  INV_X1 U2437 ( .A(n2517), .ZN(n3527) );
  AOI22_X1 U2438 ( .A1(wdata[11]), .A2(n327), .B1(n2506), .B2(x9_s1_w[11]), 
        .ZN(n2517) );
  INV_X1 U2439 ( .A(n2518), .ZN(n3511) );
  AOI22_X1 U2440 ( .A1(wdata[12]), .A2(n327), .B1(n2506), .B2(x9_s1_w[12]), 
        .ZN(n2518) );
  INV_X1 U2441 ( .A(n2519), .ZN(n3495) );
  AOI22_X1 U2442 ( .A1(wdata[13]), .A2(n327), .B1(n2506), .B2(x9_s1_w[13]), 
        .ZN(n2519) );
  INV_X1 U2443 ( .A(n2520), .ZN(n3479) );
  AOI22_X1 U2444 ( .A1(wdata[14]), .A2(n327), .B1(n2506), .B2(x9_s1_w[14]), 
        .ZN(n2520) );
  INV_X1 U2445 ( .A(n2521), .ZN(n3463) );
  AOI22_X1 U2446 ( .A1(wdata[15]), .A2(n327), .B1(n2506), .B2(x9_s1_w[15]), 
        .ZN(n2521) );
  INV_X1 U2447 ( .A(n2522), .ZN(n3447) );
  AOI22_X1 U2448 ( .A1(wdata[16]), .A2(n327), .B1(n2506), .B2(x9_s1_w[16]), 
        .ZN(n2522) );
  INV_X1 U2449 ( .A(n2523), .ZN(n3431) );
  AOI22_X1 U2450 ( .A1(wdata[17]), .A2(n327), .B1(n2506), .B2(x9_s1_w[17]), 
        .ZN(n2523) );
  INV_X1 U2451 ( .A(n2524), .ZN(n3415) );
  AOI22_X1 U2452 ( .A1(wdata[18]), .A2(n327), .B1(n2506), .B2(x9_s1_w[18]), 
        .ZN(n2524) );
  INV_X1 U2453 ( .A(n2525), .ZN(n3399) );
  AOI22_X1 U2454 ( .A1(wdata[19]), .A2(n327), .B1(n2506), .B2(x9_s1_w[19]), 
        .ZN(n2525) );
  INV_X1 U2455 ( .A(n2526), .ZN(n3383) );
  AOI22_X1 U2456 ( .A1(wdata[20]), .A2(n326), .B1(n2506), .B2(x9_s1_w[20]), 
        .ZN(n2526) );
  INV_X1 U2457 ( .A(n2527), .ZN(n3367) );
  AOI22_X1 U2458 ( .A1(wdata[21]), .A2(n326), .B1(n2506), .B2(x9_s1_w[21]), 
        .ZN(n2527) );
  INV_X1 U2459 ( .A(n2528), .ZN(n3351) );
  AOI22_X1 U2460 ( .A1(wdata[22]), .A2(n326), .B1(n2506), .B2(x9_s1_w[22]), 
        .ZN(n2528) );
  INV_X1 U2461 ( .A(n2529), .ZN(n3335) );
  AOI22_X1 U2462 ( .A1(wdata[23]), .A2(n326), .B1(n2506), .B2(x9_s1_w[23]), 
        .ZN(n2529) );
  INV_X1 U2463 ( .A(n2530), .ZN(n3319) );
  AOI22_X1 U2464 ( .A1(wdata[24]), .A2(n326), .B1(n2506), .B2(x9_s1_w[24]), 
        .ZN(n2530) );
  INV_X1 U2465 ( .A(n2531), .ZN(n3303) );
  AOI22_X1 U2466 ( .A1(wdata[25]), .A2(n326), .B1(n2506), .B2(x9_s1_w[25]), 
        .ZN(n2531) );
  INV_X1 U2467 ( .A(n2532), .ZN(n2641) );
  AOI22_X1 U2468 ( .A1(wdata[26]), .A2(n326), .B1(n2506), .B2(x9_s1_w[26]), 
        .ZN(n2532) );
  INV_X1 U2469 ( .A(n2533), .ZN(n1066) );
  AOI22_X1 U2470 ( .A1(wdata[27]), .A2(n326), .B1(n2506), .B2(x9_s1_w[27]), 
        .ZN(n2533) );
  INV_X1 U2471 ( .A(n2534), .ZN(n1050) );
  AOI22_X1 U2472 ( .A1(wdata[28]), .A2(n326), .B1(n2506), .B2(x9_s1_w[28]), 
        .ZN(n2534) );
  INV_X1 U2473 ( .A(n2535), .ZN(n1034) );
  AOI22_X1 U2474 ( .A1(wdata[29]), .A2(n326), .B1(n2506), .B2(x9_s1_w[29]), 
        .ZN(n2535) );
  INV_X1 U2475 ( .A(n2536), .ZN(n1018) );
  AOI22_X1 U2476 ( .A1(wdata[30]), .A2(n326), .B1(n2506), .B2(x9_s1_w[30]), 
        .ZN(n2536) );
  INV_X1 U2477 ( .A(n2537), .ZN(n1002) );
  AOI22_X1 U2478 ( .A1(wdata[31]), .A2(n326), .B1(n2506), .B2(x9_s1_w[31]), 
        .ZN(n2537) );
  INV_X1 U2479 ( .A(n2538), .ZN(n3702) );
  AOI22_X1 U2480 ( .A1(wdata[0]), .A2(n190), .B1(n2539), .B2(x8_s0_w[0]), .ZN(
        n2538) );
  INV_X1 U2481 ( .A(n2540), .ZN(n3686) );
  AOI22_X1 U2482 ( .A1(wdata[1]), .A2(n189), .B1(n2539), .B2(x8_s0_w[1]), .ZN(
        n2540) );
  INV_X1 U2483 ( .A(n2541), .ZN(n3670) );
  AOI22_X1 U2484 ( .A1(wdata[2]), .A2(n190), .B1(n2539), .B2(x8_s0_w[2]), .ZN(
        n2541) );
  INV_X1 U2485 ( .A(n2542), .ZN(n3654) );
  AOI22_X1 U2486 ( .A1(wdata[3]), .A2(n189), .B1(n2539), .B2(x8_s0_w[3]), .ZN(
        n2542) );
  INV_X1 U2487 ( .A(n2543), .ZN(n3638) );
  AOI22_X1 U2488 ( .A1(wdata[4]), .A2(n190), .B1(n2539), .B2(x8_s0_w[4]), .ZN(
        n2543) );
  INV_X1 U2489 ( .A(n2544), .ZN(n3622) );
  AOI22_X1 U2490 ( .A1(wdata[5]), .A2(n189), .B1(n2539), .B2(x8_s0_w[5]), .ZN(
        n2544) );
  INV_X1 U2491 ( .A(n2545), .ZN(n3606) );
  AOI22_X1 U2492 ( .A1(wdata[6]), .A2(n190), .B1(n2539), .B2(x8_s0_w[6]), .ZN(
        n2545) );
  INV_X1 U2493 ( .A(n2546), .ZN(n3590) );
  AOI22_X1 U2494 ( .A1(wdata[7]), .A2(n189), .B1(n2539), .B2(x8_s0_w[7]), .ZN(
        n2546) );
  INV_X1 U2495 ( .A(n2547), .ZN(n3574) );
  AOI22_X1 U2496 ( .A1(wdata[8]), .A2(n190), .B1(n2539), .B2(x8_s0_w[8]), .ZN(
        n2547) );
  INV_X1 U2497 ( .A(n2548), .ZN(n3558) );
  AOI22_X1 U2498 ( .A1(wdata[9]), .A2(n190), .B1(n2539), .B2(x8_s0_w[9]), .ZN(
        n2548) );
  INV_X1 U2499 ( .A(n2549), .ZN(n3542) );
  AOI22_X1 U2500 ( .A1(wdata[10]), .A2(n190), .B1(n2539), .B2(x8_s0_w[10]), 
        .ZN(n2549) );
  INV_X1 U2501 ( .A(n2550), .ZN(n3526) );
  AOI22_X1 U2502 ( .A1(wdata[11]), .A2(n190), .B1(n2539), .B2(x8_s0_w[11]), 
        .ZN(n2550) );
  INV_X1 U2503 ( .A(n2551), .ZN(n3510) );
  AOI22_X1 U2504 ( .A1(wdata[12]), .A2(n190), .B1(n2539), .B2(x8_s0_w[12]), 
        .ZN(n2551) );
  INV_X1 U2505 ( .A(n2552), .ZN(n3494) );
  AOI22_X1 U2506 ( .A1(wdata[13]), .A2(n190), .B1(n2539), .B2(x8_s0_w[13]), 
        .ZN(n2552) );
  INV_X1 U2507 ( .A(n2553), .ZN(n3478) );
  AOI22_X1 U2508 ( .A1(wdata[14]), .A2(n190), .B1(n2539), .B2(x8_s0_w[14]), 
        .ZN(n2553) );
  INV_X1 U2509 ( .A(n2554), .ZN(n3462) );
  AOI22_X1 U2510 ( .A1(wdata[15]), .A2(n190), .B1(n2539), .B2(x8_s0_w[15]), 
        .ZN(n2554) );
  INV_X1 U2511 ( .A(n2555), .ZN(n3446) );
  AOI22_X1 U2512 ( .A1(wdata[16]), .A2(n190), .B1(n2539), .B2(x8_s0_w[16]), 
        .ZN(n2555) );
  INV_X1 U2513 ( .A(n2556), .ZN(n3430) );
  AOI22_X1 U2514 ( .A1(wdata[17]), .A2(n190), .B1(n2539), .B2(x8_s0_w[17]), 
        .ZN(n2556) );
  INV_X1 U2515 ( .A(n2557), .ZN(n3414) );
  AOI22_X1 U2516 ( .A1(wdata[18]), .A2(n190), .B1(n2539), .B2(x8_s0_w[18]), 
        .ZN(n2557) );
  INV_X1 U2517 ( .A(n2558), .ZN(n3398) );
  AOI22_X1 U2518 ( .A1(wdata[19]), .A2(n190), .B1(n2539), .B2(x8_s0_w[19]), 
        .ZN(n2558) );
  INV_X1 U2519 ( .A(n2559), .ZN(n3382) );
  AOI22_X1 U2520 ( .A1(wdata[20]), .A2(n189), .B1(n2539), .B2(x8_s0_w[20]), 
        .ZN(n2559) );
  INV_X1 U2521 ( .A(n2560), .ZN(n3366) );
  AOI22_X1 U2522 ( .A1(wdata[21]), .A2(n189), .B1(n2539), .B2(x8_s0_w[21]), 
        .ZN(n2560) );
  INV_X1 U2523 ( .A(n2561), .ZN(n3350) );
  AOI22_X1 U2524 ( .A1(wdata[22]), .A2(n189), .B1(n2539), .B2(x8_s0_w[22]), 
        .ZN(n2561) );
  INV_X1 U2525 ( .A(n2562), .ZN(n3334) );
  AOI22_X1 U2526 ( .A1(wdata[23]), .A2(n189), .B1(n2539), .B2(x8_s0_w[23]), 
        .ZN(n2562) );
  INV_X1 U2527 ( .A(n2563), .ZN(n3318) );
  AOI22_X1 U2528 ( .A1(wdata[24]), .A2(n189), .B1(n2539), .B2(x8_s0_w[24]), 
        .ZN(n2563) );
  INV_X1 U2529 ( .A(n2564), .ZN(n3302) );
  AOI22_X1 U2530 ( .A1(wdata[25]), .A2(n189), .B1(n2539), .B2(x8_s0_w[25]), 
        .ZN(n2564) );
  INV_X1 U2531 ( .A(n2565), .ZN(n2640) );
  AOI22_X1 U2532 ( .A1(wdata[26]), .A2(n189), .B1(n2539), .B2(x8_s0_w[26]), 
        .ZN(n2565) );
  INV_X1 U2533 ( .A(n2566), .ZN(n1065) );
  AOI22_X1 U2534 ( .A1(wdata[27]), .A2(n189), .B1(n2539), .B2(x8_s0_w[27]), 
        .ZN(n2566) );
  INV_X1 U2535 ( .A(n2567), .ZN(n1049) );
  AOI22_X1 U2536 ( .A1(wdata[28]), .A2(n189), .B1(n2539), .B2(x8_s0_w[28]), 
        .ZN(n2567) );
  INV_X1 U2537 ( .A(n2568), .ZN(n1033) );
  AOI22_X1 U2538 ( .A1(wdata[29]), .A2(n189), .B1(n2539), .B2(x8_s0_w[29]), 
        .ZN(n2568) );
  INV_X1 U2539 ( .A(n2569), .ZN(n1017) );
  AOI22_X1 U2540 ( .A1(wdata[30]), .A2(n189), .B1(n2539), .B2(x8_s0_w[30]), 
        .ZN(n2569) );
  INV_X1 U2541 ( .A(n2570), .ZN(n1001) );
  AOI22_X1 U2542 ( .A1(wdata[31]), .A2(n189), .B1(n2539), .B2(x8_s0_w[31]), 
        .ZN(n2570) );
  INV_X1 U2543 ( .A(n2572), .ZN(n3701) );
  AOI22_X1 U2544 ( .A1(wdata[0]), .A2(n181), .B1(n2573), .B2(x7_t2_w[0]), .ZN(
        n2572) );
  INV_X1 U2545 ( .A(n2574), .ZN(n3685) );
  AOI22_X1 U2546 ( .A1(wdata[1]), .A2(n180), .B1(n2573), .B2(x7_t2_w[1]), .ZN(
        n2574) );
  INV_X1 U2547 ( .A(n2575), .ZN(n3669) );
  AOI22_X1 U2548 ( .A1(wdata[2]), .A2(n181), .B1(n2573), .B2(x7_t2_w[2]), .ZN(
        n2575) );
  INV_X1 U2549 ( .A(n2576), .ZN(n3653) );
  AOI22_X1 U2550 ( .A1(wdata[3]), .A2(n180), .B1(n2573), .B2(x7_t2_w[3]), .ZN(
        n2576) );
  INV_X1 U2551 ( .A(n2577), .ZN(n3637) );
  AOI22_X1 U2552 ( .A1(wdata[4]), .A2(n181), .B1(n2573), .B2(x7_t2_w[4]), .ZN(
        n2577) );
  INV_X1 U2553 ( .A(n2578), .ZN(n3621) );
  AOI22_X1 U2554 ( .A1(wdata[5]), .A2(n180), .B1(n2573), .B2(x7_t2_w[5]), .ZN(
        n2578) );
  INV_X1 U2555 ( .A(n2579), .ZN(n3605) );
  AOI22_X1 U2556 ( .A1(wdata[6]), .A2(n181), .B1(n2573), .B2(x7_t2_w[6]), .ZN(
        n2579) );
  INV_X1 U2557 ( .A(n2580), .ZN(n3589) );
  AOI22_X1 U2558 ( .A1(wdata[7]), .A2(n180), .B1(n2573), .B2(x7_t2_w[7]), .ZN(
        n2580) );
  INV_X1 U2559 ( .A(n2581), .ZN(n3573) );
  AOI22_X1 U2560 ( .A1(wdata[8]), .A2(n181), .B1(n2573), .B2(x7_t2_w[8]), .ZN(
        n2581) );
  INV_X1 U2561 ( .A(n2582), .ZN(n3557) );
  AOI22_X1 U2562 ( .A1(wdata[9]), .A2(n181), .B1(n2573), .B2(x7_t2_w[9]), .ZN(
        n2582) );
  INV_X1 U2563 ( .A(n2583), .ZN(n3541) );
  AOI22_X1 U2564 ( .A1(wdata[10]), .A2(n181), .B1(n2573), .B2(x7_t2_w[10]), 
        .ZN(n2583) );
  INV_X1 U2565 ( .A(n2584), .ZN(n3525) );
  AOI22_X1 U2566 ( .A1(wdata[11]), .A2(n181), .B1(n2573), .B2(x7_t2_w[11]), 
        .ZN(n2584) );
  INV_X1 U2567 ( .A(n2585), .ZN(n3509) );
  AOI22_X1 U2568 ( .A1(wdata[12]), .A2(n181), .B1(n2573), .B2(x7_t2_w[12]), 
        .ZN(n2585) );
  INV_X1 U2569 ( .A(n2586), .ZN(n3493) );
  AOI22_X1 U2570 ( .A1(wdata[13]), .A2(n181), .B1(n2573), .B2(x7_t2_w[13]), 
        .ZN(n2586) );
  INV_X1 U2571 ( .A(n2587), .ZN(n3477) );
  AOI22_X1 U2572 ( .A1(wdata[14]), .A2(n181), .B1(n2573), .B2(x7_t2_w[14]), 
        .ZN(n2587) );
  INV_X1 U2573 ( .A(n2588), .ZN(n3461) );
  AOI22_X1 U2574 ( .A1(wdata[15]), .A2(n181), .B1(n2573), .B2(x7_t2_w[15]), 
        .ZN(n2588) );
  INV_X1 U2575 ( .A(n2589), .ZN(n3445) );
  AOI22_X1 U2576 ( .A1(wdata[16]), .A2(n181), .B1(n2573), .B2(x7_t2_w[16]), 
        .ZN(n2589) );
  INV_X1 U2577 ( .A(n2590), .ZN(n3429) );
  AOI22_X1 U2578 ( .A1(wdata[17]), .A2(n181), .B1(n2573), .B2(x7_t2_w[17]), 
        .ZN(n2590) );
  INV_X1 U2579 ( .A(n2591), .ZN(n3413) );
  AOI22_X1 U2580 ( .A1(wdata[18]), .A2(n181), .B1(n2573), .B2(x7_t2_w[18]), 
        .ZN(n2591) );
  INV_X1 U2581 ( .A(n2592), .ZN(n3397) );
  AOI22_X1 U2582 ( .A1(wdata[19]), .A2(n181), .B1(n2573), .B2(x7_t2_w[19]), 
        .ZN(n2592) );
  INV_X1 U2583 ( .A(n2593), .ZN(n3381) );
  AOI22_X1 U2584 ( .A1(wdata[20]), .A2(n180), .B1(n2573), .B2(x7_t2_w[20]), 
        .ZN(n2593) );
  INV_X1 U2585 ( .A(n2594), .ZN(n3365) );
  AOI22_X1 U2586 ( .A1(wdata[21]), .A2(n180), .B1(n2573), .B2(x7_t2_w[21]), 
        .ZN(n2594) );
  INV_X1 U2587 ( .A(n2595), .ZN(n3349) );
  AOI22_X1 U2588 ( .A1(wdata[22]), .A2(n180), .B1(n2573), .B2(x7_t2_w[22]), 
        .ZN(n2595) );
  INV_X1 U2589 ( .A(n2596), .ZN(n3333) );
  AOI22_X1 U2590 ( .A1(wdata[23]), .A2(n180), .B1(n2573), .B2(x7_t2_w[23]), 
        .ZN(n2596) );
  INV_X1 U2591 ( .A(n2597), .ZN(n3317) );
  AOI22_X1 U2592 ( .A1(wdata[24]), .A2(n180), .B1(n2573), .B2(x7_t2_w[24]), 
        .ZN(n2597) );
  INV_X1 U2593 ( .A(n2598), .ZN(n3301) );
  AOI22_X1 U2594 ( .A1(wdata[25]), .A2(n180), .B1(n2573), .B2(x7_t2_w[25]), 
        .ZN(n2598) );
  INV_X1 U2595 ( .A(n2599), .ZN(n2639) );
  AOI22_X1 U2596 ( .A1(wdata[26]), .A2(n180), .B1(n2573), .B2(x7_t2_w[26]), 
        .ZN(n2599) );
  INV_X1 U2597 ( .A(n2600), .ZN(n1064) );
  AOI22_X1 U2598 ( .A1(wdata[27]), .A2(n180), .B1(n2573), .B2(x7_t2_w[27]), 
        .ZN(n2600) );
  INV_X1 U2599 ( .A(n2601), .ZN(n1048) );
  AOI22_X1 U2600 ( .A1(wdata[28]), .A2(n180), .B1(n2573), .B2(x7_t2_w[28]), 
        .ZN(n2601) );
  INV_X1 U2601 ( .A(n2602), .ZN(n1032) );
  AOI22_X1 U2602 ( .A1(wdata[29]), .A2(n180), .B1(n2573), .B2(x7_t2_w[29]), 
        .ZN(n2602) );
  INV_X1 U2603 ( .A(n2603), .ZN(n1016) );
  AOI22_X1 U2604 ( .A1(wdata[30]), .A2(n180), .B1(n2573), .B2(x7_t2_w[30]), 
        .ZN(n2603) );
  INV_X1 U2605 ( .A(n2604), .ZN(n1000) );
  AOI22_X1 U2606 ( .A1(wdata[31]), .A2(n180), .B1(n2573), .B2(x7_t2_w[31]), 
        .ZN(n2604) );
  INV_X1 U2607 ( .A(n2606), .ZN(n3700) );
  AOI22_X1 U2608 ( .A1(wdata[0]), .A2(n172), .B1(n2607), .B2(x6_t1_w[0]), .ZN(
        n2606) );
  INV_X1 U2609 ( .A(n2608), .ZN(n3684) );
  AOI22_X1 U2610 ( .A1(wdata[1]), .A2(n171), .B1(n2607), .B2(x6_t1_w[1]), .ZN(
        n2608) );
  INV_X1 U2611 ( .A(n2609), .ZN(n3668) );
  AOI22_X1 U2612 ( .A1(wdata[2]), .A2(n172), .B1(n2607), .B2(x6_t1_w[2]), .ZN(
        n2609) );
  INV_X1 U2613 ( .A(n2610), .ZN(n3652) );
  AOI22_X1 U2614 ( .A1(wdata[3]), .A2(n171), .B1(n2607), .B2(x6_t1_w[3]), .ZN(
        n2610) );
  INV_X1 U2615 ( .A(n2611), .ZN(n3636) );
  AOI22_X1 U2616 ( .A1(wdata[4]), .A2(n172), .B1(n2607), .B2(x6_t1_w[4]), .ZN(
        n2611) );
  INV_X1 U2617 ( .A(n2612), .ZN(n3620) );
  AOI22_X1 U2618 ( .A1(wdata[5]), .A2(n171), .B1(n2607), .B2(x6_t1_w[5]), .ZN(
        n2612) );
  INV_X1 U2619 ( .A(n2613), .ZN(n3604) );
  AOI22_X1 U2620 ( .A1(wdata[6]), .A2(n172), .B1(n2607), .B2(x6_t1_w[6]), .ZN(
        n2613) );
  INV_X1 U2621 ( .A(n2614), .ZN(n3588) );
  AOI22_X1 U2622 ( .A1(wdata[7]), .A2(n171), .B1(n2607), .B2(x6_t1_w[7]), .ZN(
        n2614) );
  INV_X1 U2623 ( .A(n2615), .ZN(n3572) );
  AOI22_X1 U2624 ( .A1(wdata[8]), .A2(n172), .B1(n2607), .B2(x6_t1_w[8]), .ZN(
        n2615) );
  INV_X1 U2625 ( .A(n2616), .ZN(n3556) );
  AOI22_X1 U2626 ( .A1(wdata[9]), .A2(n172), .B1(n2607), .B2(x6_t1_w[9]), .ZN(
        n2616) );
  INV_X1 U2627 ( .A(n2617), .ZN(n3540) );
  AOI22_X1 U2628 ( .A1(wdata[10]), .A2(n172), .B1(n2607), .B2(x6_t1_w[10]), 
        .ZN(n2617) );
  INV_X1 U2629 ( .A(n2618), .ZN(n3524) );
  AOI22_X1 U2630 ( .A1(wdata[11]), .A2(n172), .B1(n2607), .B2(x6_t1_w[11]), 
        .ZN(n2618) );
  INV_X1 U2631 ( .A(n2619), .ZN(n3508) );
  AOI22_X1 U2632 ( .A1(wdata[12]), .A2(n172), .B1(n2607), .B2(x6_t1_w[12]), 
        .ZN(n2619) );
  INV_X1 U2633 ( .A(n2620), .ZN(n3492) );
  AOI22_X1 U2634 ( .A1(wdata[13]), .A2(n172), .B1(n2607), .B2(x6_t1_w[13]), 
        .ZN(n2620) );
  INV_X1 U2635 ( .A(n2621), .ZN(n3476) );
  AOI22_X1 U2636 ( .A1(wdata[14]), .A2(n172), .B1(n2607), .B2(x6_t1_w[14]), 
        .ZN(n2621) );
  INV_X1 U2637 ( .A(n2622), .ZN(n3460) );
  AOI22_X1 U2638 ( .A1(wdata[15]), .A2(n172), .B1(n2607), .B2(x6_t1_w[15]), 
        .ZN(n2622) );
  INV_X1 U2639 ( .A(n2623), .ZN(n3444) );
  AOI22_X1 U2640 ( .A1(wdata[16]), .A2(n172), .B1(n2607), .B2(x6_t1_w[16]), 
        .ZN(n2623) );
  INV_X1 U2641 ( .A(n2624), .ZN(n3428) );
  AOI22_X1 U2642 ( .A1(wdata[17]), .A2(n172), .B1(n2607), .B2(x6_t1_w[17]), 
        .ZN(n2624) );
  INV_X1 U2643 ( .A(n2625), .ZN(n3412) );
  AOI22_X1 U2644 ( .A1(wdata[18]), .A2(n172), .B1(n2607), .B2(x6_t1_w[18]), 
        .ZN(n2625) );
  INV_X1 U2645 ( .A(n2626), .ZN(n3396) );
  AOI22_X1 U2646 ( .A1(wdata[19]), .A2(n172), .B1(n2607), .B2(x6_t1_w[19]), 
        .ZN(n2626) );
  INV_X1 U2647 ( .A(n2627), .ZN(n3380) );
  AOI22_X1 U2648 ( .A1(wdata[20]), .A2(n171), .B1(n2607), .B2(x6_t1_w[20]), 
        .ZN(n2627) );
  INV_X1 U2649 ( .A(n2628), .ZN(n3364) );
  AOI22_X1 U2650 ( .A1(wdata[21]), .A2(n171), .B1(n2607), .B2(x6_t1_w[21]), 
        .ZN(n2628) );
  INV_X1 U2651 ( .A(n2629), .ZN(n3348) );
  AOI22_X1 U2652 ( .A1(wdata[22]), .A2(n171), .B1(n2607), .B2(x6_t1_w[22]), 
        .ZN(n2629) );
  INV_X1 U2653 ( .A(n2630), .ZN(n3332) );
  AOI22_X1 U2654 ( .A1(wdata[23]), .A2(n171), .B1(n2607), .B2(x6_t1_w[23]), 
        .ZN(n2630) );
  INV_X1 U2655 ( .A(n2631), .ZN(n3316) );
  AOI22_X1 U2656 ( .A1(wdata[24]), .A2(n171), .B1(n2607), .B2(x6_t1_w[24]), 
        .ZN(n2631) );
  INV_X1 U2657 ( .A(n2632), .ZN(n3300) );
  AOI22_X1 U2658 ( .A1(wdata[25]), .A2(n171), .B1(n2607), .B2(x6_t1_w[25]), 
        .ZN(n2632) );
  INV_X1 U2659 ( .A(n2633), .ZN(n2504) );
  AOI22_X1 U2660 ( .A1(wdata[26]), .A2(n171), .B1(n2607), .B2(x6_t1_w[26]), 
        .ZN(n2633) );
  INV_X1 U2661 ( .A(n2634), .ZN(n1063) );
  AOI22_X1 U2662 ( .A1(wdata[27]), .A2(n171), .B1(n2607), .B2(x6_t1_w[27]), 
        .ZN(n2634) );
  INV_X1 U2663 ( .A(n2635), .ZN(n1047) );
  AOI22_X1 U2664 ( .A1(wdata[28]), .A2(n171), .B1(n2607), .B2(x6_t1_w[28]), 
        .ZN(n2635) );
  INV_X1 U2665 ( .A(n2636), .ZN(n1031) );
  AOI22_X1 U2666 ( .A1(wdata[29]), .A2(n171), .B1(n2607), .B2(x6_t1_w[29]), 
        .ZN(n2636) );
  INV_X1 U2667 ( .A(n2637), .ZN(n1015) );
  AOI22_X1 U2668 ( .A1(wdata[30]), .A2(n171), .B1(n2607), .B2(x6_t1_w[30]), 
        .ZN(n2637) );
  INV_X1 U2669 ( .A(n2638), .ZN(n999) );
  AOI22_X1 U2670 ( .A1(wdata[31]), .A2(n171), .B1(n2607), .B2(x6_t1_w[31]), 
        .ZN(n2638) );
  INV_X1 U2671 ( .A(n2644), .ZN(n3699) );
  AOI22_X1 U2672 ( .A1(wdata[0]), .A2(n127), .B1(n2645), .B2(x1_ra_w[0]), .ZN(
        n2644) );
  INV_X1 U2673 ( .A(n2646), .ZN(n3683) );
  AOI22_X1 U2674 ( .A1(wdata[1]), .A2(n126), .B1(n2645), .B2(x1_ra_w[1]), .ZN(
        n2646) );
  INV_X1 U2675 ( .A(n2647), .ZN(n3667) );
  AOI22_X1 U2676 ( .A1(wdata[2]), .A2(n127), .B1(n2645), .B2(x1_ra_w[2]), .ZN(
        n2647) );
  INV_X1 U2677 ( .A(n2648), .ZN(n3651) );
  AOI22_X1 U2678 ( .A1(wdata[3]), .A2(n126), .B1(n2645), .B2(x1_ra_w[3]), .ZN(
        n2648) );
  INV_X1 U2679 ( .A(n2649), .ZN(n3635) );
  AOI22_X1 U2680 ( .A1(wdata[4]), .A2(n127), .B1(n2645), .B2(x1_ra_w[4]), .ZN(
        n2649) );
  INV_X1 U2681 ( .A(n2650), .ZN(n3619) );
  AOI22_X1 U2682 ( .A1(wdata[5]), .A2(n126), .B1(n2645), .B2(x1_ra_w[5]), .ZN(
        n2650) );
  INV_X1 U2683 ( .A(n2651), .ZN(n3603) );
  AOI22_X1 U2684 ( .A1(wdata[6]), .A2(n127), .B1(n2645), .B2(x1_ra_w[6]), .ZN(
        n2651) );
  INV_X1 U2685 ( .A(n2652), .ZN(n3587) );
  AOI22_X1 U2686 ( .A1(wdata[7]), .A2(n126), .B1(n2645), .B2(x1_ra_w[7]), .ZN(
        n2652) );
  INV_X1 U2687 ( .A(n2653), .ZN(n3571) );
  AOI22_X1 U2688 ( .A1(wdata[8]), .A2(n127), .B1(n2645), .B2(x1_ra_w[8]), .ZN(
        n2653) );
  INV_X1 U2689 ( .A(n2654), .ZN(n3555) );
  AOI22_X1 U2690 ( .A1(wdata[9]), .A2(n127), .B1(n2645), .B2(x1_ra_w[9]), .ZN(
        n2654) );
  INV_X1 U2691 ( .A(n2655), .ZN(n3539) );
  AOI22_X1 U2692 ( .A1(wdata[10]), .A2(n127), .B1(n2645), .B2(x1_ra_w[10]), 
        .ZN(n2655) );
  INV_X1 U2693 ( .A(n2656), .ZN(n3523) );
  AOI22_X1 U2694 ( .A1(wdata[11]), .A2(n127), .B1(n2645), .B2(x1_ra_w[11]), 
        .ZN(n2656) );
  INV_X1 U2695 ( .A(n2657), .ZN(n3507) );
  AOI22_X1 U2696 ( .A1(wdata[12]), .A2(n127), .B1(n2645), .B2(x1_ra_w[12]), 
        .ZN(n2657) );
  INV_X1 U2697 ( .A(n2658), .ZN(n3491) );
  AOI22_X1 U2698 ( .A1(wdata[13]), .A2(n127), .B1(n2645), .B2(x1_ra_w[13]), 
        .ZN(n2658) );
  INV_X1 U2699 ( .A(n2659), .ZN(n3475) );
  AOI22_X1 U2700 ( .A1(wdata[14]), .A2(n127), .B1(n2645), .B2(x1_ra_w[14]), 
        .ZN(n2659) );
  INV_X1 U2701 ( .A(n2660), .ZN(n3459) );
  AOI22_X1 U2702 ( .A1(wdata[15]), .A2(n127), .B1(n2645), .B2(x1_ra_w[15]), 
        .ZN(n2660) );
  INV_X1 U2703 ( .A(n2661), .ZN(n3443) );
  AOI22_X1 U2704 ( .A1(wdata[16]), .A2(n127), .B1(n2645), .B2(x1_ra_w[16]), 
        .ZN(n2661) );
  INV_X1 U2705 ( .A(n2662), .ZN(n3427) );
  AOI22_X1 U2706 ( .A1(wdata[17]), .A2(n127), .B1(n2645), .B2(x1_ra_w[17]), 
        .ZN(n2662) );
  INV_X1 U2707 ( .A(n2663), .ZN(n3411) );
  AOI22_X1 U2708 ( .A1(wdata[18]), .A2(n127), .B1(n2645), .B2(x1_ra_w[18]), 
        .ZN(n2663) );
  INV_X1 U2709 ( .A(n2664), .ZN(n3395) );
  AOI22_X1 U2710 ( .A1(wdata[19]), .A2(n127), .B1(n2645), .B2(x1_ra_w[19]), 
        .ZN(n2664) );
  INV_X1 U2711 ( .A(n2665), .ZN(n3379) );
  AOI22_X1 U2712 ( .A1(wdata[20]), .A2(n126), .B1(n2645), .B2(x1_ra_w[20]), 
        .ZN(n2665) );
  INV_X1 U2713 ( .A(n2666), .ZN(n3363) );
  AOI22_X1 U2714 ( .A1(wdata[21]), .A2(n126), .B1(n2645), .B2(x1_ra_w[21]), 
        .ZN(n2666) );
  INV_X1 U2715 ( .A(n2667), .ZN(n3347) );
  AOI22_X1 U2716 ( .A1(wdata[22]), .A2(n126), .B1(n2645), .B2(x1_ra_w[22]), 
        .ZN(n2667) );
  INV_X1 U2717 ( .A(n2668), .ZN(n3331) );
  AOI22_X1 U2718 ( .A1(wdata[23]), .A2(n126), .B1(n2645), .B2(x1_ra_w[23]), 
        .ZN(n2668) );
  INV_X1 U2719 ( .A(n2669), .ZN(n3315) );
  AOI22_X1 U2720 ( .A1(wdata[24]), .A2(n126), .B1(n2645), .B2(x1_ra_w[24]), 
        .ZN(n2669) );
  INV_X1 U2721 ( .A(n2670), .ZN(n3299) );
  AOI22_X1 U2722 ( .A1(wdata[25]), .A2(n126), .B1(n2645), .B2(x1_ra_w[25]), 
        .ZN(n2670) );
  INV_X1 U2723 ( .A(n2671), .ZN(n2502) );
  AOI22_X1 U2724 ( .A1(wdata[26]), .A2(n126), .B1(n2645), .B2(x1_ra_w[26]), 
        .ZN(n2671) );
  INV_X1 U2725 ( .A(n2672), .ZN(n1062) );
  AOI22_X1 U2726 ( .A1(wdata[27]), .A2(n126), .B1(n2645), .B2(x1_ra_w[27]), 
        .ZN(n2672) );
  INV_X1 U2727 ( .A(n2673), .ZN(n1046) );
  AOI22_X1 U2728 ( .A1(wdata[28]), .A2(n126), .B1(n2645), .B2(x1_ra_w[28]), 
        .ZN(n2673) );
  INV_X1 U2729 ( .A(n2674), .ZN(n1030) );
  AOI22_X1 U2730 ( .A1(wdata[29]), .A2(n126), .B1(n2645), .B2(x1_ra_w[29]), 
        .ZN(n2674) );
  INV_X1 U2731 ( .A(n2675), .ZN(n1014) );
  AOI22_X1 U2732 ( .A1(wdata[30]), .A2(n126), .B1(n2645), .B2(x1_ra_w[30]), 
        .ZN(n2675) );
  INV_X1 U2733 ( .A(n2676), .ZN(n998) );
  AOI22_X1 U2734 ( .A1(wdata[31]), .A2(n126), .B1(n2645), .B2(x1_ra_w[31]), 
        .ZN(n2676) );
  INV_X1 U2735 ( .A(n2677), .ZN(n3698) );
  AOI22_X1 U2736 ( .A1(wdata[0]), .A2(n118), .B1(n2678), .B2(x31_t6_w[0]), 
        .ZN(n2677) );
  INV_X1 U2737 ( .A(n2679), .ZN(n3682) );
  AOI22_X1 U2738 ( .A1(wdata[1]), .A2(n117), .B1(n2678), .B2(x31_t6_w[1]), 
        .ZN(n2679) );
  INV_X1 U2739 ( .A(n2680), .ZN(n3666) );
  AOI22_X1 U2740 ( .A1(wdata[2]), .A2(n118), .B1(n2678), .B2(x31_t6_w[2]), 
        .ZN(n2680) );
  INV_X1 U2741 ( .A(n2681), .ZN(n3650) );
  AOI22_X1 U2742 ( .A1(wdata[3]), .A2(n117), .B1(n2678), .B2(x31_t6_w[3]), 
        .ZN(n2681) );
  INV_X1 U2743 ( .A(n2682), .ZN(n3634) );
  AOI22_X1 U2744 ( .A1(wdata[4]), .A2(n118), .B1(n2678), .B2(x31_t6_w[4]), 
        .ZN(n2682) );
  INV_X1 U2745 ( .A(n2683), .ZN(n3618) );
  AOI22_X1 U2746 ( .A1(wdata[5]), .A2(n117), .B1(n2678), .B2(x31_t6_w[5]), 
        .ZN(n2683) );
  INV_X1 U2747 ( .A(n2684), .ZN(n3602) );
  AOI22_X1 U2748 ( .A1(wdata[6]), .A2(n118), .B1(n2678), .B2(x31_t6_w[6]), 
        .ZN(n2684) );
  INV_X1 U2749 ( .A(n2685), .ZN(n3586) );
  AOI22_X1 U2750 ( .A1(wdata[7]), .A2(n117), .B1(n2678), .B2(x31_t6_w[7]), 
        .ZN(n2685) );
  INV_X1 U2751 ( .A(n2686), .ZN(n3570) );
  AOI22_X1 U2752 ( .A1(wdata[8]), .A2(n118), .B1(n2678), .B2(x31_t6_w[8]), 
        .ZN(n2686) );
  INV_X1 U2753 ( .A(n2687), .ZN(n3554) );
  AOI22_X1 U2754 ( .A1(wdata[9]), .A2(n118), .B1(n2678), .B2(x31_t6_w[9]), 
        .ZN(n2687) );
  INV_X1 U2755 ( .A(n2688), .ZN(n3538) );
  AOI22_X1 U2756 ( .A1(wdata[10]), .A2(n118), .B1(n2678), .B2(x31_t6_w[10]), 
        .ZN(n2688) );
  INV_X1 U2757 ( .A(n2689), .ZN(n3522) );
  AOI22_X1 U2758 ( .A1(wdata[11]), .A2(n118), .B1(n2678), .B2(x31_t6_w[11]), 
        .ZN(n2689) );
  INV_X1 U2759 ( .A(n2690), .ZN(n3506) );
  AOI22_X1 U2760 ( .A1(wdata[12]), .A2(n118), .B1(n2678), .B2(x31_t6_w[12]), 
        .ZN(n2690) );
  INV_X1 U2761 ( .A(n2691), .ZN(n3490) );
  AOI22_X1 U2762 ( .A1(wdata[13]), .A2(n118), .B1(n2678), .B2(x31_t6_w[13]), 
        .ZN(n2691) );
  INV_X1 U2763 ( .A(n2692), .ZN(n3474) );
  AOI22_X1 U2764 ( .A1(wdata[14]), .A2(n118), .B1(n2678), .B2(x31_t6_w[14]), 
        .ZN(n2692) );
  INV_X1 U2765 ( .A(n2693), .ZN(n3458) );
  AOI22_X1 U2766 ( .A1(wdata[15]), .A2(n118), .B1(n2678), .B2(x31_t6_w[15]), 
        .ZN(n2693) );
  INV_X1 U2767 ( .A(n2694), .ZN(n3442) );
  AOI22_X1 U2768 ( .A1(wdata[16]), .A2(n118), .B1(n2678), .B2(x31_t6_w[16]), 
        .ZN(n2694) );
  INV_X1 U2769 ( .A(n2695), .ZN(n3426) );
  AOI22_X1 U2770 ( .A1(wdata[17]), .A2(n118), .B1(n2678), .B2(x31_t6_w[17]), 
        .ZN(n2695) );
  INV_X1 U2771 ( .A(n2696), .ZN(n3410) );
  AOI22_X1 U2772 ( .A1(wdata[18]), .A2(n118), .B1(n2678), .B2(x31_t6_w[18]), 
        .ZN(n2696) );
  INV_X1 U2773 ( .A(n2697), .ZN(n3394) );
  AOI22_X1 U2774 ( .A1(wdata[19]), .A2(n118), .B1(n2678), .B2(x31_t6_w[19]), 
        .ZN(n2697) );
  INV_X1 U2775 ( .A(n2698), .ZN(n3378) );
  AOI22_X1 U2776 ( .A1(wdata[20]), .A2(n117), .B1(n2678), .B2(x31_t6_w[20]), 
        .ZN(n2698) );
  INV_X1 U2777 ( .A(n2699), .ZN(n3362) );
  AOI22_X1 U2778 ( .A1(wdata[21]), .A2(n117), .B1(n2678), .B2(x31_t6_w[21]), 
        .ZN(n2699) );
  INV_X1 U2779 ( .A(n2700), .ZN(n3346) );
  AOI22_X1 U2844 ( .A1(wdata[22]), .A2(n117), .B1(n2678), .B2(x31_t6_w[22]), 
        .ZN(n2700) );
  INV_X1 U2845 ( .A(n2701), .ZN(n3330) );
  AOI22_X1 U2846 ( .A1(wdata[23]), .A2(n117), .B1(n2678), .B2(x31_t6_w[23]), 
        .ZN(n2701) );
  INV_X1 U2847 ( .A(n2702), .ZN(n3314) );
  AOI22_X1 U2848 ( .A1(wdata[24]), .A2(n117), .B1(n2678), .B2(x31_t6_w[24]), 
        .ZN(n2702) );
  INV_X1 U2849 ( .A(n2703), .ZN(n3298) );
  AOI22_X1 U2850 ( .A1(wdata[25]), .A2(n117), .B1(n2678), .B2(x31_t6_w[25]), 
        .ZN(n2703) );
  INV_X1 U2851 ( .A(n2704), .ZN(n2499) );
  AOI22_X1 U2852 ( .A1(wdata[26]), .A2(n117), .B1(n2678), .B2(x31_t6_w[26]), 
        .ZN(n2704) );
  INV_X1 U2853 ( .A(n2705), .ZN(n1061) );
  AOI22_X1 U2854 ( .A1(wdata[27]), .A2(n117), .B1(n2678), .B2(x31_t6_w[27]), 
        .ZN(n2705) );
  INV_X1 U2855 ( .A(n2706), .ZN(n1045) );
  AOI22_X1 U2856 ( .A1(wdata[28]), .A2(n117), .B1(n2678), .B2(x31_t6_w[28]), 
        .ZN(n2706) );
  INV_X1 U2857 ( .A(n2707), .ZN(n1029) );
  AOI22_X1 U2858 ( .A1(wdata[29]), .A2(n117), .B1(n2678), .B2(x31_t6_w[29]), 
        .ZN(n2707) );
  INV_X1 U2859 ( .A(n2708), .ZN(n1013) );
  AOI22_X1 U2860 ( .A1(wdata[30]), .A2(n117), .B1(n2678), .B2(x31_t6_w[30]), 
        .ZN(n2708) );
  INV_X1 U2861 ( .A(n2709), .ZN(n997) );
  AOI22_X1 U2862 ( .A1(wdata[31]), .A2(n117), .B1(n2678), .B2(x31_t6_w[31]), 
        .ZN(n2709) );
  INV_X1 U2863 ( .A(n2711), .ZN(n3697) );
  AOI22_X1 U2864 ( .A1(wdata[0]), .A2(n109), .B1(n2712), .B2(x30_t5_w[0]), 
        .ZN(n2711) );
  INV_X1 U2865 ( .A(n2713), .ZN(n3681) );
  AOI22_X1 U2866 ( .A1(wdata[1]), .A2(n108), .B1(n2712), .B2(x30_t5_w[1]), 
        .ZN(n2713) );
  INV_X1 U2867 ( .A(n2714), .ZN(n3665) );
  AOI22_X1 U2868 ( .A1(wdata[2]), .A2(n109), .B1(n2712), .B2(x30_t5_w[2]), 
        .ZN(n2714) );
  INV_X1 U2869 ( .A(n2715), .ZN(n3649) );
  AOI22_X1 U2870 ( .A1(wdata[3]), .A2(n108), .B1(n2712), .B2(x30_t5_w[3]), 
        .ZN(n2715) );
  INV_X1 U2871 ( .A(n2716), .ZN(n3633) );
  AOI22_X1 U2872 ( .A1(wdata[4]), .A2(n109), .B1(n2712), .B2(x30_t5_w[4]), 
        .ZN(n2716) );
  INV_X1 U2873 ( .A(n2717), .ZN(n3617) );
  AOI22_X1 U2874 ( .A1(wdata[5]), .A2(n108), .B1(n2712), .B2(x30_t5_w[5]), 
        .ZN(n2717) );
  INV_X1 U2875 ( .A(n2718), .ZN(n3601) );
  AOI22_X1 U2876 ( .A1(wdata[6]), .A2(n109), .B1(n2712), .B2(x30_t5_w[6]), 
        .ZN(n2718) );
  INV_X1 U2877 ( .A(n2719), .ZN(n3585) );
  AOI22_X1 U2878 ( .A1(wdata[7]), .A2(n108), .B1(n2712), .B2(x30_t5_w[7]), 
        .ZN(n2719) );
  INV_X1 U2879 ( .A(n2720), .ZN(n3569) );
  AOI22_X1 U2880 ( .A1(wdata[8]), .A2(n109), .B1(n2712), .B2(x30_t5_w[8]), 
        .ZN(n2720) );
  INV_X1 U2881 ( .A(n2721), .ZN(n3553) );
  AOI22_X1 U2882 ( .A1(wdata[9]), .A2(n109), .B1(n2712), .B2(x30_t5_w[9]), 
        .ZN(n2721) );
  INV_X1 U2883 ( .A(n2722), .ZN(n3537) );
  AOI22_X1 U2884 ( .A1(wdata[10]), .A2(n109), .B1(n2712), .B2(x30_t5_w[10]), 
        .ZN(n2722) );
  INV_X1 U2885 ( .A(n2723), .ZN(n3521) );
  AOI22_X1 U2886 ( .A1(wdata[11]), .A2(n109), .B1(n2712), .B2(x30_t5_w[11]), 
        .ZN(n2723) );
  INV_X1 U2887 ( .A(n2724), .ZN(n3505) );
  AOI22_X1 U2888 ( .A1(wdata[12]), .A2(n109), .B1(n2712), .B2(x30_t5_w[12]), 
        .ZN(n2724) );
  INV_X1 U2889 ( .A(n2725), .ZN(n3489) );
  AOI22_X1 U2890 ( .A1(wdata[13]), .A2(n109), .B1(n2712), .B2(x30_t5_w[13]), 
        .ZN(n2725) );
  INV_X1 U2891 ( .A(n2726), .ZN(n3473) );
  AOI22_X1 U2892 ( .A1(wdata[14]), .A2(n109), .B1(n2712), .B2(x30_t5_w[14]), 
        .ZN(n2726) );
  INV_X1 U2893 ( .A(n2727), .ZN(n3457) );
  AOI22_X1 U2894 ( .A1(wdata[15]), .A2(n109), .B1(n2712), .B2(x30_t5_w[15]), 
        .ZN(n2727) );
  INV_X1 U2895 ( .A(n2728), .ZN(n3441) );
  AOI22_X1 U2896 ( .A1(wdata[16]), .A2(n109), .B1(n2712), .B2(x30_t5_w[16]), 
        .ZN(n2728) );
  INV_X1 U2897 ( .A(n2729), .ZN(n3425) );
  AOI22_X1 U2898 ( .A1(wdata[17]), .A2(n109), .B1(n2712), .B2(x30_t5_w[17]), 
        .ZN(n2729) );
  INV_X1 U2899 ( .A(n2730), .ZN(n3409) );
  AOI22_X1 U2900 ( .A1(wdata[18]), .A2(n109), .B1(n2712), .B2(x30_t5_w[18]), 
        .ZN(n2730) );
  INV_X1 U2901 ( .A(n2731), .ZN(n3393) );
  AOI22_X1 U2902 ( .A1(wdata[19]), .A2(n109), .B1(n2712), .B2(x30_t5_w[19]), 
        .ZN(n2731) );
  INV_X1 U2903 ( .A(n2732), .ZN(n3377) );
  AOI22_X1 U2904 ( .A1(wdata[20]), .A2(n108), .B1(n2712), .B2(x30_t5_w[20]), 
        .ZN(n2732) );
  INV_X1 U2905 ( .A(n2733), .ZN(n3361) );
  AOI22_X1 U2906 ( .A1(wdata[21]), .A2(n108), .B1(n2712), .B2(x30_t5_w[21]), 
        .ZN(n2733) );
  INV_X1 U2907 ( .A(n2734), .ZN(n3345) );
  AOI22_X1 U2908 ( .A1(wdata[22]), .A2(n108), .B1(n2712), .B2(x30_t5_w[22]), 
        .ZN(n2734) );
  INV_X1 U2909 ( .A(n2735), .ZN(n3329) );
  AOI22_X1 U2910 ( .A1(wdata[23]), .A2(n108), .B1(n2712), .B2(x30_t5_w[23]), 
        .ZN(n2735) );
  INV_X1 U2911 ( .A(n2736), .ZN(n3313) );
  AOI22_X1 U2912 ( .A1(wdata[24]), .A2(n108), .B1(n2712), .B2(x30_t5_w[24]), 
        .ZN(n2736) );
  INV_X1 U2913 ( .A(n2737), .ZN(n3297) );
  AOI22_X1 U2914 ( .A1(wdata[25]), .A2(n108), .B1(n2712), .B2(x30_t5_w[25]), 
        .ZN(n2737) );
  INV_X1 U2915 ( .A(n2738), .ZN(n2498) );
  AOI22_X1 U2916 ( .A1(wdata[26]), .A2(n108), .B1(n2712), .B2(x30_t5_w[26]), 
        .ZN(n2738) );
  INV_X1 U2917 ( .A(n2739), .ZN(n1060) );
  AOI22_X1 U2918 ( .A1(wdata[27]), .A2(n108), .B1(n2712), .B2(x30_t5_w[27]), 
        .ZN(n2739) );
  INV_X1 U2919 ( .A(n2740), .ZN(n1044) );
  AOI22_X1 U2920 ( .A1(wdata[28]), .A2(n108), .B1(n2712), .B2(x30_t5_w[28]), 
        .ZN(n2740) );
  INV_X1 U2921 ( .A(n2741), .ZN(n1028) );
  AOI22_X1 U2922 ( .A1(wdata[29]), .A2(n108), .B1(n2712), .B2(x30_t5_w[29]), 
        .ZN(n2741) );
  INV_X1 U2923 ( .A(n2742), .ZN(n1012) );
  AOI22_X1 U2924 ( .A1(wdata[30]), .A2(n108), .B1(n2712), .B2(x30_t5_w[30]), 
        .ZN(n2742) );
  INV_X1 U2925 ( .A(n2743), .ZN(n996) );
  AOI22_X1 U2926 ( .A1(wdata[31]), .A2(n108), .B1(n2712), .B2(x30_t5_w[31]), 
        .ZN(n2743) );
  INV_X1 U2927 ( .A(n2744), .ZN(n3696) );
  AOI22_X1 U2928 ( .A1(wdata[0]), .A2(n100), .B1(n2745), .B2(x27_s11_w[0]), 
        .ZN(n2744) );
  INV_X1 U2929 ( .A(n2746), .ZN(n3680) );
  AOI22_X1 U2930 ( .A1(wdata[1]), .A2(n99), .B1(n2745), .B2(x27_s11_w[1]), 
        .ZN(n2746) );
  INV_X1 U2931 ( .A(n2747), .ZN(n3664) );
  AOI22_X1 U2932 ( .A1(wdata[2]), .A2(n100), .B1(n2745), .B2(x27_s11_w[2]), 
        .ZN(n2747) );
  INV_X1 U2933 ( .A(n2748), .ZN(n3648) );
  AOI22_X1 U2934 ( .A1(wdata[3]), .A2(n99), .B1(n2745), .B2(x27_s11_w[3]), 
        .ZN(n2748) );
  INV_X1 U2935 ( .A(n2749), .ZN(n3632) );
  AOI22_X1 U2936 ( .A1(wdata[4]), .A2(n100), .B1(n2745), .B2(x27_s11_w[4]), 
        .ZN(n2749) );
  INV_X1 U2937 ( .A(n2750), .ZN(n3616) );
  AOI22_X1 U2938 ( .A1(wdata[5]), .A2(n99), .B1(n2745), .B2(x27_s11_w[5]), 
        .ZN(n2750) );
  INV_X1 U2939 ( .A(n2751), .ZN(n3600) );
  AOI22_X1 U2940 ( .A1(wdata[6]), .A2(n100), .B1(n2745), .B2(x27_s11_w[6]), 
        .ZN(n2751) );
  INV_X1 U2941 ( .A(n2752), .ZN(n3584) );
  AOI22_X1 U2942 ( .A1(wdata[7]), .A2(n99), .B1(n2745), .B2(x27_s11_w[7]), 
        .ZN(n2752) );
  INV_X1 U2943 ( .A(n2753), .ZN(n3568) );
  AOI22_X1 U2944 ( .A1(wdata[8]), .A2(n100), .B1(n2745), .B2(x27_s11_w[8]), 
        .ZN(n2753) );
  INV_X1 U2945 ( .A(n2754), .ZN(n3552) );
  AOI22_X1 U2946 ( .A1(wdata[9]), .A2(n100), .B1(n2745), .B2(x27_s11_w[9]), 
        .ZN(n2754) );
  INV_X1 U2947 ( .A(n2755), .ZN(n3536) );
  AOI22_X1 U2948 ( .A1(wdata[10]), .A2(n100), .B1(n2745), .B2(x27_s11_w[10]), 
        .ZN(n2755) );
  INV_X1 U2949 ( .A(n2756), .ZN(n3520) );
  AOI22_X1 U2950 ( .A1(wdata[11]), .A2(n100), .B1(n2745), .B2(x27_s11_w[11]), 
        .ZN(n2756) );
  INV_X1 U2951 ( .A(n2757), .ZN(n3504) );
  AOI22_X1 U2952 ( .A1(wdata[12]), .A2(n100), .B1(n2745), .B2(x27_s11_w[12]), 
        .ZN(n2757) );
  INV_X1 U2953 ( .A(n2758), .ZN(n3488) );
  AOI22_X1 U2954 ( .A1(wdata[13]), .A2(n100), .B1(n2745), .B2(x27_s11_w[13]), 
        .ZN(n2758) );
  INV_X1 U2955 ( .A(n2759), .ZN(n3472) );
  AOI22_X1 U2956 ( .A1(wdata[14]), .A2(n100), .B1(n2745), .B2(x27_s11_w[14]), 
        .ZN(n2759) );
  INV_X1 U2957 ( .A(n2760), .ZN(n3456) );
  AOI22_X1 U2958 ( .A1(wdata[15]), .A2(n100), .B1(n2745), .B2(x27_s11_w[15]), 
        .ZN(n2760) );
  INV_X1 U2959 ( .A(n2761), .ZN(n3440) );
  AOI22_X1 U2960 ( .A1(wdata[16]), .A2(n100), .B1(n2745), .B2(x27_s11_w[16]), 
        .ZN(n2761) );
  INV_X1 U2961 ( .A(n2762), .ZN(n3424) );
  AOI22_X1 U2962 ( .A1(wdata[17]), .A2(n100), .B1(n2745), .B2(x27_s11_w[17]), 
        .ZN(n2762) );
  INV_X1 U2963 ( .A(n2763), .ZN(n3408) );
  AOI22_X1 U2964 ( .A1(wdata[18]), .A2(n100), .B1(n2745), .B2(x27_s11_w[18]), 
        .ZN(n2763) );
  INV_X1 U2965 ( .A(n2764), .ZN(n3392) );
  AOI22_X1 U2966 ( .A1(wdata[19]), .A2(n100), .B1(n2745), .B2(x27_s11_w[19]), 
        .ZN(n2764) );
  INV_X1 U2967 ( .A(n2765), .ZN(n3376) );
  AOI22_X1 U2968 ( .A1(wdata[20]), .A2(n99), .B1(n2745), .B2(x27_s11_w[20]), 
        .ZN(n2765) );
  INV_X1 U2969 ( .A(n2766), .ZN(n3360) );
  AOI22_X1 U2970 ( .A1(wdata[21]), .A2(n99), .B1(n2745), .B2(x27_s11_w[21]), 
        .ZN(n2766) );
  INV_X1 U2971 ( .A(n2767), .ZN(n3344) );
  AOI22_X1 U2972 ( .A1(wdata[22]), .A2(n99), .B1(n2745), .B2(x27_s11_w[22]), 
        .ZN(n2767) );
  INV_X1 U2973 ( .A(n2768), .ZN(n3328) );
  AOI22_X1 U2974 ( .A1(wdata[23]), .A2(n99), .B1(n2745), .B2(x27_s11_w[23]), 
        .ZN(n2768) );
  INV_X1 U2975 ( .A(n2769), .ZN(n3312) );
  AOI22_X1 U2976 ( .A1(wdata[24]), .A2(n99), .B1(n2745), .B2(x27_s11_w[24]), 
        .ZN(n2769) );
  INV_X1 U2977 ( .A(n2770), .ZN(n3296) );
  AOI22_X1 U2978 ( .A1(wdata[25]), .A2(n99), .B1(n2745), .B2(x27_s11_w[25]), 
        .ZN(n2770) );
  INV_X1 U2979 ( .A(n2771), .ZN(n2363) );
  AOI22_X1 U2980 ( .A1(wdata[26]), .A2(n99), .B1(n2745), .B2(x27_s11_w[26]), 
        .ZN(n2771) );
  INV_X1 U2981 ( .A(n2772), .ZN(n1059) );
  AOI22_X1 U2982 ( .A1(wdata[27]), .A2(n99), .B1(n2745), .B2(x27_s11_w[27]), 
        .ZN(n2772) );
  INV_X1 U2983 ( .A(n2773), .ZN(n1043) );
  AOI22_X1 U2984 ( .A1(wdata[28]), .A2(n99), .B1(n2745), .B2(x27_s11_w[28]), 
        .ZN(n2773) );
  INV_X1 U2985 ( .A(n2774), .ZN(n1027) );
  AOI22_X1 U2986 ( .A1(wdata[29]), .A2(n99), .B1(n2745), .B2(x27_s11_w[29]), 
        .ZN(n2774) );
  INV_X1 U2987 ( .A(n2775), .ZN(n1011) );
  AOI22_X1 U2988 ( .A1(wdata[30]), .A2(n99), .B1(n2745), .B2(x27_s11_w[30]), 
        .ZN(n2775) );
  INV_X1 U2989 ( .A(n2776), .ZN(n995) );
  AOI22_X1 U2990 ( .A1(wdata[31]), .A2(n99), .B1(n2745), .B2(x27_s11_w[31]), 
        .ZN(n2776) );
  INV_X1 U2991 ( .A(n2250), .ZN(n3710) );
  AOI22_X1 U2992 ( .A1(n608), .A2(wdata[0]), .B1(n2251), .B2(x26_s10_w[0]), 
        .ZN(n2250) );
  INV_X1 U2993 ( .A(n2252), .ZN(n3694) );
  AOI22_X1 U2994 ( .A1(n607), .A2(wdata[1]), .B1(n2251), .B2(x26_s10_w[1]), 
        .ZN(n2252) );
  INV_X1 U2995 ( .A(n2253), .ZN(n3678) );
  AOI22_X1 U2996 ( .A1(n608), .A2(wdata[2]), .B1(n2251), .B2(x26_s10_w[2]), 
        .ZN(n2253) );
  INV_X1 U2997 ( .A(n2254), .ZN(n3662) );
  AOI22_X1 U2998 ( .A1(n607), .A2(wdata[3]), .B1(n2251), .B2(x26_s10_w[3]), 
        .ZN(n2254) );
  INV_X1 U2999 ( .A(n2255), .ZN(n3646) );
  AOI22_X1 U3000 ( .A1(n608), .A2(wdata[4]), .B1(n2251), .B2(x26_s10_w[4]), 
        .ZN(n2255) );
  INV_X1 U3001 ( .A(n2256), .ZN(n3630) );
  AOI22_X1 U3002 ( .A1(n607), .A2(wdata[5]), .B1(n2251), .B2(x26_s10_w[5]), 
        .ZN(n2256) );
  INV_X1 U3003 ( .A(n2257), .ZN(n3614) );
  AOI22_X1 U3004 ( .A1(n608), .A2(wdata[6]), .B1(n2251), .B2(x26_s10_w[6]), 
        .ZN(n2257) );
  INV_X1 U3005 ( .A(n2258), .ZN(n3598) );
  AOI22_X1 U3006 ( .A1(n607), .A2(wdata[7]), .B1(n2251), .B2(x26_s10_w[7]), 
        .ZN(n2258) );
  INV_X1 U3007 ( .A(n2259), .ZN(n3582) );
  AOI22_X1 U3008 ( .A1(n608), .A2(wdata[8]), .B1(n2251), .B2(x26_s10_w[8]), 
        .ZN(n2259) );
  INV_X1 U3009 ( .A(n2260), .ZN(n3566) );
  AOI22_X1 U3010 ( .A1(n608), .A2(wdata[9]), .B1(n2251), .B2(x26_s10_w[9]), 
        .ZN(n2260) );
  INV_X1 U3011 ( .A(n2261), .ZN(n3550) );
  AOI22_X1 U3012 ( .A1(n608), .A2(wdata[10]), .B1(n2251), .B2(x26_s10_w[10]), 
        .ZN(n2261) );
  INV_X1 U3013 ( .A(n2262), .ZN(n3534) );
  AOI22_X1 U3014 ( .A1(n608), .A2(wdata[11]), .B1(n2251), .B2(x26_s10_w[11]), 
        .ZN(n2262) );
  INV_X1 U3015 ( .A(n2263), .ZN(n3518) );
  AOI22_X1 U3016 ( .A1(n608), .A2(wdata[12]), .B1(n2251), .B2(x26_s10_w[12]), 
        .ZN(n2263) );
  INV_X1 U3017 ( .A(n2264), .ZN(n3502) );
  AOI22_X1 U3018 ( .A1(n608), .A2(wdata[13]), .B1(n2251), .B2(x26_s10_w[13]), 
        .ZN(n2264) );
  INV_X1 U3019 ( .A(n2265), .ZN(n3486) );
  AOI22_X1 U3020 ( .A1(n608), .A2(wdata[14]), .B1(n2251), .B2(x26_s10_w[14]), 
        .ZN(n2265) );
  INV_X1 U3021 ( .A(n2266), .ZN(n3470) );
  AOI22_X1 U3022 ( .A1(n608), .A2(wdata[15]), .B1(n2251), .B2(x26_s10_w[15]), 
        .ZN(n2266) );
  INV_X1 U3023 ( .A(n2267), .ZN(n3454) );
  AOI22_X1 U3024 ( .A1(n608), .A2(wdata[16]), .B1(n2251), .B2(x26_s10_w[16]), 
        .ZN(n2267) );
  INV_X1 U3025 ( .A(n2268), .ZN(n3438) );
  AOI22_X1 U3026 ( .A1(n608), .A2(wdata[17]), .B1(n2251), .B2(x26_s10_w[17]), 
        .ZN(n2268) );
  INV_X1 U3027 ( .A(n2269), .ZN(n3422) );
  AOI22_X1 U3028 ( .A1(n608), .A2(wdata[18]), .B1(n2251), .B2(x26_s10_w[18]), 
        .ZN(n2269) );
  INV_X1 U3029 ( .A(n2270), .ZN(n3406) );
  AOI22_X1 U3030 ( .A1(n608), .A2(wdata[19]), .B1(n2251), .B2(x26_s10_w[19]), 
        .ZN(n2270) );
  INV_X1 U3031 ( .A(n2271), .ZN(n3390) );
  AOI22_X1 U3032 ( .A1(n607), .A2(wdata[20]), .B1(n2251), .B2(x26_s10_w[20]), 
        .ZN(n2271) );
  INV_X1 U3033 ( .A(n2272), .ZN(n3374) );
  AOI22_X1 U3034 ( .A1(n607), .A2(wdata[21]), .B1(n2251), .B2(x26_s10_w[21]), 
        .ZN(n2272) );
  INV_X1 U3035 ( .A(n2273), .ZN(n3358) );
  AOI22_X1 U3036 ( .A1(n607), .A2(wdata[22]), .B1(n2251), .B2(x26_s10_w[22]), 
        .ZN(n2273) );
  INV_X1 U3037 ( .A(n2274), .ZN(n3342) );
  AOI22_X1 U3038 ( .A1(n607), .A2(wdata[23]), .B1(n2251), .B2(x26_s10_w[23]), 
        .ZN(n2274) );
  INV_X1 U3039 ( .A(n2275), .ZN(n3326) );
  AOI22_X1 U3040 ( .A1(n607), .A2(wdata[24]), .B1(n2251), .B2(x26_s10_w[24]), 
        .ZN(n2275) );
  INV_X1 U3041 ( .A(n2276), .ZN(n3310) );
  AOI22_X1 U3042 ( .A1(n607), .A2(wdata[25]), .B1(n2251), .B2(x26_s10_w[25]), 
        .ZN(n2276) );
  INV_X1 U3043 ( .A(n2277), .ZN(n3294) );
  AOI22_X1 U3044 ( .A1(n607), .A2(wdata[26]), .B1(n2251), .B2(x26_s10_w[26]), 
        .ZN(n2277) );
  INV_X1 U3045 ( .A(n2278), .ZN(n2358) );
  AOI22_X1 U3046 ( .A1(n607), .A2(wdata[27]), .B1(n2251), .B2(x26_s10_w[27]), 
        .ZN(n2278) );
  INV_X1 U3047 ( .A(n2279), .ZN(n1057) );
  AOI22_X1 U3048 ( .A1(n607), .A2(wdata[28]), .B1(n2251), .B2(x26_s10_w[28]), 
        .ZN(n2279) );
  INV_X1 U3049 ( .A(n2280), .ZN(n1041) );
  AOI22_X1 U3050 ( .A1(n607), .A2(wdata[29]), .B1(n2251), .B2(x26_s10_w[29]), 
        .ZN(n2280) );
  INV_X1 U3051 ( .A(n2281), .ZN(n1025) );
  AOI22_X1 U3052 ( .A1(n607), .A2(wdata[30]), .B1(n2251), .B2(x26_s10_w[30]), 
        .ZN(n2281) );
  INV_X1 U3053 ( .A(n2282), .ZN(n1009) );
  AOI22_X1 U3054 ( .A1(n607), .A2(wdata[31]), .B1(n2251), .B2(x26_s10_w[31]), 
        .ZN(n2282) );
  OAI22_X1 U3055 ( .A1(n1111), .A2(n544), .B1(n1112), .B2(n576), .ZN(n1657) );
  OAI22_X1 U3056 ( .A1(n1116), .A2(n480), .B1(n1117), .B2(n512), .ZN(n1658) );
  OAI22_X1 U3057 ( .A1(n1111), .A2(n543), .B1(n1112), .B2(n575), .ZN(n1456) );
  OAI22_X1 U3058 ( .A1(n1116), .A2(n479), .B1(n1117), .B2(n511), .ZN(n1457) );
  OAI22_X1 U3059 ( .A1(n1111), .A2(n542), .B1(n1112), .B2(n574), .ZN(n1269) );
  OAI22_X1 U3060 ( .A1(n1116), .A2(n478), .B1(n1117), .B2(n510), .ZN(n1270) );
  OAI22_X1 U3061 ( .A1(n1111), .A2(n534), .B1(n1112), .B2(n566), .ZN(n1626) );
  OAI22_X1 U3062 ( .A1(n1116), .A2(n470), .B1(n1117), .B2(n502), .ZN(n1627) );
  OAI22_X1 U3063 ( .A1(n1111), .A2(n533), .B1(n1112), .B2(n565), .ZN(n1609) );
  OAI22_X1 U3064 ( .A1(n1116), .A2(n469), .B1(n1117), .B2(n501), .ZN(n1610) );
  OAI22_X1 U3065 ( .A1(n1111), .A2(n532), .B1(n1112), .B2(n564), .ZN(n1592) );
  OAI22_X1 U3066 ( .A1(n1116), .A2(n468), .B1(n1117), .B2(n500), .ZN(n1593) );
  OAI22_X1 U3067 ( .A1(n1111), .A2(n531), .B1(n1112), .B2(n563), .ZN(n1575) );
  OAI22_X1 U3068 ( .A1(n1116), .A2(n467), .B1(n1117), .B2(n499), .ZN(n1576) );
  OAI22_X1 U3069 ( .A1(n1111), .A2(n530), .B1(n1112), .B2(n562), .ZN(n1558) );
  OAI22_X1 U3070 ( .A1(n1116), .A2(n466), .B1(n1117), .B2(n498), .ZN(n1559) );
  OAI22_X1 U3071 ( .A1(n1111), .A2(n529), .B1(n1112), .B2(n561), .ZN(n1541) );
  OAI22_X1 U3072 ( .A1(n1116), .A2(n465), .B1(n1117), .B2(n497), .ZN(n1542) );
  OAI22_X1 U3073 ( .A1(n1111), .A2(n528), .B1(n1112), .B2(n560), .ZN(n1524) );
  OAI22_X1 U3074 ( .A1(n1116), .A2(n464), .B1(n1117), .B2(n496), .ZN(n1525) );
  OAI22_X1 U3075 ( .A1(n1111), .A2(n527), .B1(n1112), .B2(n559), .ZN(n1507) );
  OAI22_X1 U3076 ( .A1(n1116), .A2(n463), .B1(n1117), .B2(n495), .ZN(n1508) );
  OAI22_X1 U3077 ( .A1(n1111), .A2(n526), .B1(n1112), .B2(n558), .ZN(n1490) );
  OAI22_X1 U3078 ( .A1(n1116), .A2(n462), .B1(n1117), .B2(n494), .ZN(n1491) );
  OAI22_X1 U3079 ( .A1(n1111), .A2(n525), .B1(n1112), .B2(n557), .ZN(n1473) );
  OAI22_X1 U3080 ( .A1(n1116), .A2(n461), .B1(n1117), .B2(n493), .ZN(n1474) );
  OAI22_X1 U3081 ( .A1(n1111), .A2(n524), .B1(n1112), .B2(n556), .ZN(n1439) );
  OAI22_X1 U3082 ( .A1(n1116), .A2(n460), .B1(n1117), .B2(n492), .ZN(n1440) );
  OAI22_X1 U3083 ( .A1(n1111), .A2(n523), .B1(n1112), .B2(n555), .ZN(n1422) );
  OAI22_X1 U3084 ( .A1(n1116), .A2(n459), .B1(n1117), .B2(n491), .ZN(n1423) );
  OAI22_X1 U3085 ( .A1(n1111), .A2(n522), .B1(n1112), .B2(n554), .ZN(n1405) );
  OAI22_X1 U3086 ( .A1(n1116), .A2(n458), .B1(n1117), .B2(n490), .ZN(n1406) );
  OAI22_X1 U3087 ( .A1(n1111), .A2(n521), .B1(n1112), .B2(n553), .ZN(n1388) );
  OAI22_X1 U3088 ( .A1(n1116), .A2(n457), .B1(n1117), .B2(n489), .ZN(n1389) );
  OAI22_X1 U3089 ( .A1(n1111), .A2(n520), .B1(n1112), .B2(n552), .ZN(n1371) );
  OAI22_X1 U3090 ( .A1(n1116), .A2(n456), .B1(n1117), .B2(n488), .ZN(n1372) );
  OAI22_X1 U3091 ( .A1(n1111), .A2(n519), .B1(n1112), .B2(n551), .ZN(n1354) );
  OAI22_X1 U3092 ( .A1(n1116), .A2(n455), .B1(n1117), .B2(n487), .ZN(n1355) );
  OAI22_X1 U3093 ( .A1(n1111), .A2(n518), .B1(n1112), .B2(n550), .ZN(n1337) );
  OAI22_X1 U3094 ( .A1(n1116), .A2(n454), .B1(n1117), .B2(n486), .ZN(n1338) );
  OAI22_X1 U3095 ( .A1(n1111), .A2(n517), .B1(n1112), .B2(n549), .ZN(n1320) );
  OAI22_X1 U3096 ( .A1(n1116), .A2(n453), .B1(n1117), .B2(n485), .ZN(n1321) );
  OAI22_X1 U3097 ( .A1(n1111), .A2(n516), .B1(n1112), .B2(n548), .ZN(n1303) );
  OAI22_X1 U3098 ( .A1(n1116), .A2(n452), .B1(n1117), .B2(n484), .ZN(n1304) );
  OAI22_X1 U3099 ( .A1(n1111), .A2(n515), .B1(n1112), .B2(n547), .ZN(n1286) );
  OAI22_X1 U3100 ( .A1(n1116), .A2(n451), .B1(n1117), .B2(n483), .ZN(n1287) );
  OAI22_X1 U3101 ( .A1(n1111), .A2(n514), .B1(n1112), .B2(n546), .ZN(n1252) );
  OAI22_X1 U3102 ( .A1(n1116), .A2(n450), .B1(n1117), .B2(n482), .ZN(n1253) );
  OAI22_X1 U3103 ( .A1(n544), .A2(n1701), .B1(n576), .B2(n1702), .ZN(n2247) );
  OAI22_X1 U3104 ( .A1(n480), .A2(n1706), .B1(n512), .B2(n1707), .ZN(n2248) );
  OAI22_X1 U3105 ( .A1(n543), .A2(n1701), .B1(n575), .B2(n1702), .ZN(n2046) );
  OAI22_X1 U3106 ( .A1(n479), .A2(n1706), .B1(n511), .B2(n1707), .ZN(n2047) );
  OAI22_X1 U3107 ( .A1(n542), .A2(n1701), .B1(n574), .B2(n1702), .ZN(n1859) );
  OAI22_X1 U3108 ( .A1(n478), .A2(n1706), .B1(n510), .B2(n1707), .ZN(n1860) );
  OAI22_X1 U3109 ( .A1(n541), .A2(n1701), .B1(n573), .B2(n1702), .ZN(n1808) );
  OAI22_X1 U3110 ( .A1(n477), .A2(n1706), .B1(n509), .B2(n1707), .ZN(n1809) );
  OAI22_X1 U3111 ( .A1(n540), .A2(n1701), .B1(n572), .B2(n1702), .ZN(n1791) );
  OAI22_X1 U3112 ( .A1(n476), .A2(n1706), .B1(n508), .B2(n1707), .ZN(n1792) );
  OAI22_X1 U3113 ( .A1(n539), .A2(n1701), .B1(n571), .B2(n1702), .ZN(n1774) );
  OAI22_X1 U3114 ( .A1(n475), .A2(n1706), .B1(n507), .B2(n1707), .ZN(n1775) );
  OAI22_X1 U3115 ( .A1(n538), .A2(n1701), .B1(n570), .B2(n1702), .ZN(n1757) );
  OAI22_X1 U3116 ( .A1(n474), .A2(n1706), .B1(n506), .B2(n1707), .ZN(n1758) );
  OAI22_X1 U3117 ( .A1(n537), .A2(n1701), .B1(n569), .B2(n1702), .ZN(n1740) );
  OAI22_X1 U3118 ( .A1(n473), .A2(n1706), .B1(n505), .B2(n1707), .ZN(n1741) );
  OAI22_X1 U3119 ( .A1(n536), .A2(n1701), .B1(n568), .B2(n1702), .ZN(n1723) );
  OAI22_X1 U3120 ( .A1(n472), .A2(n1706), .B1(n504), .B2(n1707), .ZN(n1724) );
  OAI22_X1 U3121 ( .A1(n535), .A2(n1701), .B1(n567), .B2(n1702), .ZN(n1700) );
  OAI22_X1 U3122 ( .A1(n471), .A2(n1706), .B1(n503), .B2(n1707), .ZN(n1705) );
  OAI22_X1 U3123 ( .A1(n534), .A2(n1701), .B1(n566), .B2(n1702), .ZN(n2216) );
  OAI22_X1 U3124 ( .A1(n470), .A2(n1706), .B1(n502), .B2(n1707), .ZN(n2217) );
  OAI22_X1 U3125 ( .A1(n533), .A2(n1701), .B1(n565), .B2(n1702), .ZN(n2199) );
  OAI22_X1 U3126 ( .A1(n469), .A2(n1706), .B1(n501), .B2(n1707), .ZN(n2200) );
  OAI22_X1 U3127 ( .A1(n532), .A2(n1701), .B1(n564), .B2(n1702), .ZN(n2182) );
  OAI22_X1 U3128 ( .A1(n468), .A2(n1706), .B1(n500), .B2(n1707), .ZN(n2183) );
  OAI22_X1 U3129 ( .A1(n531), .A2(n1701), .B1(n563), .B2(n1702), .ZN(n2165) );
  OAI22_X1 U3130 ( .A1(n467), .A2(n1706), .B1(n499), .B2(n1707), .ZN(n2166) );
  OAI22_X1 U3131 ( .A1(n530), .A2(n1701), .B1(n562), .B2(n1702), .ZN(n2148) );
  OAI22_X1 U3132 ( .A1(n466), .A2(n1706), .B1(n498), .B2(n1707), .ZN(n2149) );
  OAI22_X1 U3133 ( .A1(n529), .A2(n1701), .B1(n561), .B2(n1702), .ZN(n2131) );
  OAI22_X1 U3134 ( .A1(n465), .A2(n1706), .B1(n497), .B2(n1707), .ZN(n2132) );
  OAI22_X1 U3135 ( .A1(n528), .A2(n1701), .B1(n560), .B2(n1702), .ZN(n2114) );
  OAI22_X1 U3136 ( .A1(n464), .A2(n1706), .B1(n496), .B2(n1707), .ZN(n2115) );
  OAI22_X1 U3137 ( .A1(n527), .A2(n1701), .B1(n559), .B2(n1702), .ZN(n2097) );
  OAI22_X1 U3138 ( .A1(n463), .A2(n1706), .B1(n495), .B2(n1707), .ZN(n2098) );
  OAI22_X1 U3139 ( .A1(n526), .A2(n1701), .B1(n558), .B2(n1702), .ZN(n2080) );
  OAI22_X1 U3140 ( .A1(n462), .A2(n1706), .B1(n494), .B2(n1707), .ZN(n2081) );
  OAI22_X1 U3141 ( .A1(n525), .A2(n1701), .B1(n557), .B2(n1702), .ZN(n2063) );
  OAI22_X1 U3142 ( .A1(n461), .A2(n1706), .B1(n493), .B2(n1707), .ZN(n2064) );
  OAI22_X1 U3143 ( .A1(n524), .A2(n1701), .B1(n556), .B2(n1702), .ZN(n2029) );
  OAI22_X1 U3144 ( .A1(n460), .A2(n1706), .B1(n492), .B2(n1707), .ZN(n2030) );
  OAI22_X1 U3145 ( .A1(n523), .A2(n1701), .B1(n555), .B2(n1702), .ZN(n2012) );
  OAI22_X1 U3146 ( .A1(n459), .A2(n1706), .B1(n491), .B2(n1707), .ZN(n2013) );
  OAI22_X1 U3147 ( .A1(n522), .A2(n1701), .B1(n554), .B2(n1702), .ZN(n1995) );
  OAI22_X1 U3148 ( .A1(n458), .A2(n1706), .B1(n490), .B2(n1707), .ZN(n1996) );
  OAI22_X1 U3149 ( .A1(n521), .A2(n1701), .B1(n553), .B2(n1702), .ZN(n1978) );
  OAI22_X1 U3150 ( .A1(n457), .A2(n1706), .B1(n489), .B2(n1707), .ZN(n1979) );
  OAI22_X1 U3151 ( .A1(n520), .A2(n1701), .B1(n552), .B2(n1702), .ZN(n1961) );
  OAI22_X1 U3152 ( .A1(n456), .A2(n1706), .B1(n488), .B2(n1707), .ZN(n1962) );
  OAI22_X1 U3153 ( .A1(n519), .A2(n1701), .B1(n551), .B2(n1702), .ZN(n1944) );
  OAI22_X1 U3154 ( .A1(n455), .A2(n1706), .B1(n487), .B2(n1707), .ZN(n1945) );
  OAI22_X1 U3155 ( .A1(n518), .A2(n1701), .B1(n550), .B2(n1702), .ZN(n1927) );
  OAI22_X1 U3156 ( .A1(n454), .A2(n1706), .B1(n486), .B2(n1707), .ZN(n1928) );
  OAI22_X1 U3157 ( .A1(n517), .A2(n1701), .B1(n549), .B2(n1702), .ZN(n1910) );
  OAI22_X1 U3158 ( .A1(n453), .A2(n1706), .B1(n485), .B2(n1707), .ZN(n1911) );
  OAI22_X1 U3159 ( .A1(n516), .A2(n1701), .B1(n548), .B2(n1702), .ZN(n1893) );
  OAI22_X1 U3160 ( .A1(n452), .A2(n1706), .B1(n484), .B2(n1707), .ZN(n1894) );
  OAI22_X1 U3161 ( .A1(n515), .A2(n1701), .B1(n547), .B2(n1702), .ZN(n1876) );
  OAI22_X1 U3162 ( .A1(n451), .A2(n1706), .B1(n483), .B2(n1707), .ZN(n1877) );
  OAI22_X1 U3163 ( .A1(n514), .A2(n1701), .B1(n546), .B2(n1702), .ZN(n1842) );
  OAI22_X1 U3164 ( .A1(n450), .A2(n1706), .B1(n482), .B2(n1707), .ZN(n1843) );
  OAI22_X1 U3165 ( .A1(n513), .A2(n1701), .B1(n545), .B2(n1702), .ZN(n1825) );
  OAI22_X1 U3166 ( .A1(n449), .A2(n1706), .B1(n481), .B2(n1707), .ZN(n1826) );
  OAI22_X1 U3167 ( .A1(n1111), .A2(n541), .B1(n1112), .B2(n573), .ZN(n1218) );
  OAI22_X1 U3168 ( .A1(n1116), .A2(n477), .B1(n1117), .B2(n509), .ZN(n1219) );
  OAI22_X1 U3169 ( .A1(n1111), .A2(n540), .B1(n1112), .B2(n572), .ZN(n1201) );
  OAI22_X1 U3170 ( .A1(n1116), .A2(n476), .B1(n1117), .B2(n508), .ZN(n1202) );
  OAI22_X1 U3171 ( .A1(n1111), .A2(n539), .B1(n1112), .B2(n571), .ZN(n1184) );
  OAI22_X1 U3172 ( .A1(n1116), .A2(n475), .B1(n1117), .B2(n507), .ZN(n1185) );
  OAI22_X1 U3173 ( .A1(n1111), .A2(n538), .B1(n1112), .B2(n570), .ZN(n1167) );
  OAI22_X1 U3174 ( .A1(n1116), .A2(n474), .B1(n1117), .B2(n506), .ZN(n1168) );
  OAI22_X1 U3175 ( .A1(n1111), .A2(n537), .B1(n1112), .B2(n569), .ZN(n1150) );
  OAI22_X1 U3176 ( .A1(n1116), .A2(n473), .B1(n1117), .B2(n505), .ZN(n1151) );
  OAI22_X1 U3177 ( .A1(n1111), .A2(n536), .B1(n1112), .B2(n568), .ZN(n1133) );
  OAI22_X1 U3178 ( .A1(n1116), .A2(n472), .B1(n1117), .B2(n504), .ZN(n1134) );
  OAI22_X1 U3179 ( .A1(n1111), .A2(n535), .B1(n1112), .B2(n567), .ZN(n1110) );
  OAI22_X1 U3180 ( .A1(n1116), .A2(n471), .B1(n1117), .B2(n503), .ZN(n1115) );
  OAI22_X1 U3181 ( .A1(n1111), .A2(n513), .B1(n1112), .B2(n545), .ZN(n1235) );
  OAI22_X1 U3182 ( .A1(n1116), .A2(n449), .B1(n1117), .B2(n481), .ZN(n1236) );
  OAI22_X1 U3183 ( .A1(n1101), .A2(n224), .B1(n1102), .B2(n256), .ZN(n1651) );
  OAI22_X1 U3184 ( .A1(n1101), .A2(n223), .B1(n1102), .B2(n255), .ZN(n1454) );
  OAI22_X1 U3185 ( .A1(n1101), .A2(n222), .B1(n1102), .B2(n254), .ZN(n1267) );
  OAI22_X1 U3186 ( .A1(n1101), .A2(n214), .B1(n1102), .B2(n246), .ZN(n1624) );
  OAI22_X1 U3187 ( .A1(n1101), .A2(n213), .B1(n1102), .B2(n245), .ZN(n1607) );
  OAI22_X1 U3188 ( .A1(n1101), .A2(n212), .B1(n1102), .B2(n244), .ZN(n1590) );
  OAI22_X1 U3189 ( .A1(n1101), .A2(n211), .B1(n1102), .B2(n243), .ZN(n1573) );
  OAI22_X1 U3190 ( .A1(n1101), .A2(n210), .B1(n1102), .B2(n242), .ZN(n1556) );
  OAI22_X1 U3191 ( .A1(n1101), .A2(n209), .B1(n1102), .B2(n241), .ZN(n1539) );
  OAI22_X1 U3192 ( .A1(n1101), .A2(n208), .B1(n1102), .B2(n240), .ZN(n1522) );
  OAI22_X1 U3193 ( .A1(n1101), .A2(n207), .B1(n1102), .B2(n239), .ZN(n1505) );
  OAI22_X1 U3194 ( .A1(n1101), .A2(n206), .B1(n1102), .B2(n238), .ZN(n1488) );
  OAI22_X1 U3195 ( .A1(n1101), .A2(n205), .B1(n1102), .B2(n237), .ZN(n1471) );
  OAI22_X1 U3196 ( .A1(n1101), .A2(n204), .B1(n1102), .B2(n236), .ZN(n1437) );
  OAI22_X1 U3197 ( .A1(n1101), .A2(n203), .B1(n1102), .B2(n235), .ZN(n1420) );
  OAI22_X1 U3198 ( .A1(n1101), .A2(n202), .B1(n1102), .B2(n234), .ZN(n1403) );
  OAI22_X1 U3199 ( .A1(n1101), .A2(n201), .B1(n1102), .B2(n233), .ZN(n1386) );
  OAI22_X1 U3200 ( .A1(n1101), .A2(n200), .B1(n1102), .B2(n232), .ZN(n1369) );
  OAI22_X1 U3201 ( .A1(n1101), .A2(n199), .B1(n1102), .B2(n231), .ZN(n1352) );
  OAI22_X1 U3202 ( .A1(n1101), .A2(n198), .B1(n1102), .B2(n230), .ZN(n1335) );
  OAI22_X1 U3203 ( .A1(n1101), .A2(n197), .B1(n1102), .B2(n229), .ZN(n1318) );
  OAI22_X1 U3204 ( .A1(n1101), .A2(n196), .B1(n1102), .B2(n228), .ZN(n1301) );
  OAI22_X1 U3205 ( .A1(n1101), .A2(n195), .B1(n1102), .B2(n227), .ZN(n1284) );
  OAI22_X1 U3206 ( .A1(n1101), .A2(n194), .B1(n1102), .B2(n226), .ZN(n1250) );
  OAI22_X1 U3207 ( .A1(n224), .A2(n1691), .B1(n256), .B2(n1692), .ZN(n2241) );
  OAI22_X1 U3208 ( .A1(n223), .A2(n1691), .B1(n255), .B2(n1692), .ZN(n2044) );
  OAI22_X1 U3209 ( .A1(n222), .A2(n1691), .B1(n254), .B2(n1692), .ZN(n1857) );
  OAI22_X1 U3210 ( .A1(n221), .A2(n1691), .B1(n253), .B2(n1692), .ZN(n1806) );
  OAI22_X1 U3211 ( .A1(n220), .A2(n1691), .B1(n252), .B2(n1692), .ZN(n1789) );
  OAI22_X1 U3212 ( .A1(n219), .A2(n1691), .B1(n251), .B2(n1692), .ZN(n1772) );
  OAI22_X1 U3213 ( .A1(n218), .A2(n1691), .B1(n250), .B2(n1692), .ZN(n1755) );
  OAI22_X1 U3214 ( .A1(n217), .A2(n1691), .B1(n249), .B2(n1692), .ZN(n1738) );
  OAI22_X1 U3215 ( .A1(n216), .A2(n1691), .B1(n248), .B2(n1692), .ZN(n1721) );
  OAI22_X1 U3216 ( .A1(n215), .A2(n1691), .B1(n247), .B2(n1692), .ZN(n1690) );
  OAI22_X1 U3217 ( .A1(n214), .A2(n1691), .B1(n246), .B2(n1692), .ZN(n2214) );
  OAI22_X1 U3218 ( .A1(n213), .A2(n1691), .B1(n245), .B2(n1692), .ZN(n2197) );
  OAI22_X1 U3219 ( .A1(n212), .A2(n1691), .B1(n244), .B2(n1692), .ZN(n2180) );
  OAI22_X1 U3220 ( .A1(n211), .A2(n1691), .B1(n243), .B2(n1692), .ZN(n2163) );
  OAI22_X1 U3221 ( .A1(n210), .A2(n1691), .B1(n242), .B2(n1692), .ZN(n2146) );
  OAI22_X1 U3222 ( .A1(n209), .A2(n1691), .B1(n241), .B2(n1692), .ZN(n2129) );
  OAI22_X1 U3223 ( .A1(n208), .A2(n1691), .B1(n240), .B2(n1692), .ZN(n2112) );
  OAI22_X1 U3224 ( .A1(n207), .A2(n1691), .B1(n239), .B2(n1692), .ZN(n2095) );
  OAI22_X1 U3225 ( .A1(n206), .A2(n1691), .B1(n238), .B2(n1692), .ZN(n2078) );
  OAI22_X1 U3226 ( .A1(n205), .A2(n1691), .B1(n237), .B2(n1692), .ZN(n2061) );
  OAI22_X1 U3227 ( .A1(n204), .A2(n1691), .B1(n236), .B2(n1692), .ZN(n2027) );
  OAI22_X1 U3228 ( .A1(n203), .A2(n1691), .B1(n235), .B2(n1692), .ZN(n2010) );
  OAI22_X1 U3229 ( .A1(n202), .A2(n1691), .B1(n234), .B2(n1692), .ZN(n1993) );
  OAI22_X1 U3230 ( .A1(n201), .A2(n1691), .B1(n233), .B2(n1692), .ZN(n1976) );
  OAI22_X1 U3231 ( .A1(n200), .A2(n1691), .B1(n232), .B2(n1692), .ZN(n1959) );
  OAI22_X1 U3232 ( .A1(n199), .A2(n1691), .B1(n231), .B2(n1692), .ZN(n1942) );
  OAI22_X1 U3233 ( .A1(n198), .A2(n1691), .B1(n230), .B2(n1692), .ZN(n1925) );
  OAI22_X1 U3234 ( .A1(n197), .A2(n1691), .B1(n229), .B2(n1692), .ZN(n1908) );
  OAI22_X1 U3235 ( .A1(n196), .A2(n1691), .B1(n228), .B2(n1692), .ZN(n1891) );
  OAI22_X1 U3236 ( .A1(n195), .A2(n1691), .B1(n227), .B2(n1692), .ZN(n1874) );
  OAI22_X1 U3237 ( .A1(n194), .A2(n1691), .B1(n226), .B2(n1692), .ZN(n1840) );
  OAI22_X1 U3238 ( .A1(n193), .A2(n1691), .B1(n225), .B2(n1692), .ZN(n1823) );
  OAI22_X1 U3239 ( .A1(n1101), .A2(n221), .B1(n1102), .B2(n253), .ZN(n1216) );
  OAI22_X1 U3240 ( .A1(n1101), .A2(n220), .B1(n1102), .B2(n252), .ZN(n1199) );
  OAI22_X1 U3241 ( .A1(n1101), .A2(n219), .B1(n1102), .B2(n251), .ZN(n1182) );
  OAI22_X1 U3242 ( .A1(n1101), .A2(n218), .B1(n1102), .B2(n250), .ZN(n1165) );
  OAI22_X1 U3243 ( .A1(n1101), .A2(n217), .B1(n1102), .B2(n249), .ZN(n1148) );
  OAI22_X1 U3244 ( .A1(n1101), .A2(n216), .B1(n1102), .B2(n248), .ZN(n1131) );
  OAI22_X1 U3245 ( .A1(n1101), .A2(n215), .B1(n1102), .B2(n247), .ZN(n1100) );
  OAI22_X1 U3246 ( .A1(n1101), .A2(n193), .B1(n1102), .B2(n225), .ZN(n1233) );
  NOR2_X1 U3247 ( .A1(n3719), .A2(ra2[4]), .ZN(n1652) );
  NOR2_X1 U3248 ( .A1(n3723), .A2(ra1[4]), .ZN(n2242) );
  NOR2_X1 U3249 ( .A1(ra2[4]), .A2(ra2[0]), .ZN(n1653) );
  NOR2_X1 U3250 ( .A1(ra1[4]), .A2(ra1[0]), .ZN(n2243) );
  NOR3_X1 U3251 ( .A1(ra2[2]), .A2(ra2[3]), .A3(ra2[1]), .ZN(n1637) );
  NOR3_X1 U3252 ( .A1(ra1[2]), .A2(ra1[3]), .A3(ra1[1]), .ZN(n2227) );
  AND2_X1 U3253 ( .A1(ra2[4]), .A2(ra2[0]), .ZN(n1639) );
  AND2_X1 U3254 ( .A1(ra1[4]), .A2(ra1[0]), .ZN(n2229) );
  AND2_X1 U3255 ( .A1(ra2[4]), .A2(n3719), .ZN(n1638) );
  AND2_X1 U3256 ( .A1(ra1[4]), .A2(n3723), .ZN(n2228) );
  AND2_X1 U3257 ( .A1(n1656), .A2(ra2[3]), .ZN(n1649) );
  AND2_X1 U3258 ( .A1(n2246), .A2(ra1[3]), .ZN(n2239) );
  NOR2_X1 U3259 ( .A1(n3717), .A2(ra2[1]), .ZN(n1656) );
  NOR2_X1 U3260 ( .A1(n3721), .A2(ra1[1]), .ZN(n2246) );
  NOR2_X1 U3261 ( .A1(n3718), .A2(ra2[3]), .ZN(n1654) );
  NOR2_X1 U3262 ( .A1(n3722), .A2(ra1[3]), .ZN(n2244) );
  NOR2_X1 U3263 ( .A1(n3716), .A2(ra2[2]), .ZN(n1659) );
  NOR2_X1 U3264 ( .A1(n3720), .A2(ra1[2]), .ZN(n2249) );
  AND2_X1 U3265 ( .A1(n1659), .A2(ra2[1]), .ZN(n1645) );
  AND2_X1 U3266 ( .A1(n2249), .A2(ra1[1]), .ZN(n2235) );
  INV_X1 U3267 ( .A(ra2[3]), .ZN(n3716) );
  INV_X1 U3268 ( .A(ra1[3]), .ZN(n3720) );
  INV_X1 U3269 ( .A(ra2[1]), .ZN(n3718) );
  INV_X1 U3270 ( .A(ra1[1]), .ZN(n3722) );
  INV_X1 U3271 ( .A(ra2[2]), .ZN(n3717) );
  INV_X1 U3272 ( .A(ra1[2]), .ZN(n3721) );
  AND2_X1 U3273 ( .A1(n1654), .A2(ra2[2]), .ZN(n1642) );
  AND2_X1 U3274 ( .A1(n2244), .A2(ra1[2]), .ZN(n2232) );
  INV_X1 U3275 ( .A(ra2[0]), .ZN(n3719) );
  INV_X1 U3276 ( .A(ra1[0]), .ZN(n3723) );
  INV_X2 U3277 ( .A(clk), .ZN(n3724) );
  INV_X2 U16 ( .A(n82), .ZN(n80) );
  NAND2_X1 U18 ( .A1(n2710), .A2(n2288), .ZN(n82) );
  INV_X2 U20 ( .A(n154), .ZN(n68) );
  NAND2_X1 U40 ( .A1(n2605), .A2(n2288), .ZN(n154) );
  INV_X2 U42 ( .A(n354), .ZN(n79) );
  NAND2_X1 U44 ( .A1(n2464), .A2(n2288), .ZN(n354) );
  INV_X2 U46 ( .A(n426), .ZN(n78) );
  NAND2_X1 U48 ( .A1(n2323), .A2(n2288), .ZN(n426) );
  INV_X2 U50 ( .A(n590), .ZN(n69) );
  NAND2_X1 U52 ( .A1(n2288), .A2(n2284), .ZN(n590) );
  INV_X2 U54 ( .A(n91), .ZN(n77) );
  NAND2_X1 U56 ( .A1(n2710), .A2(n2286), .ZN(n91) );
  INV_X2 U58 ( .A(n163), .ZN(n75) );
  NAND2_X1 U60 ( .A1(n2605), .A2(n2286), .ZN(n163) );
  INV_X2 U62 ( .A(n363), .ZN(n73) );
  NAND2_X1 U64 ( .A1(n2464), .A2(n2286), .ZN(n363) );
  INV_X2 U68 ( .A(n435), .ZN(n71) );
  NAND2_X1 U69 ( .A1(n2323), .A2(n2286), .ZN(n435) );
  INV_X2 U70 ( .A(n136), .ZN(n76) );
  NAND2_X1 U71 ( .A1(n2642), .A2(n2283), .ZN(n136) );
  INV_X2 U72 ( .A(n599), .ZN(n70) );
  NAND2_X1 U73 ( .A1(n2286), .A2(n2284), .ZN(n599) );
  INV_X2 U74 ( .A(n145), .ZN(n67) );
  NAND2_X1 U75 ( .A1(n2642), .A2(n2322), .ZN(n145) );
  INV_X2 U76 ( .A(n336), .ZN(n74) );
  NAND2_X1 U77 ( .A1(n2503), .A2(n2283), .ZN(n336) );
  INV_X2 U78 ( .A(n408), .ZN(n72) );
  NAND2_X1 U79 ( .A1(n2362), .A2(n2283), .ZN(n408) );
  INV_X2 U80 ( .A(n345), .ZN(n66) );
  NAND2_X1 U81 ( .A1(n2503), .A2(n2322), .ZN(n345) );
  INV_X2 U82 ( .A(n417), .ZN(n65) );
  NAND2_X1 U83 ( .A1(n2362), .A2(n2322), .ZN(n417) );
  NAND2_X2 U84 ( .A1(n2284), .A2(n2322), .ZN(n2745) );
  NAND2_X2 U85 ( .A1(n2323), .A2(n2322), .ZN(n2290) );
  NAND2_X2 U86 ( .A1(n2288), .A2(n2503), .ZN(n2539) );
  NAND2_X2 U87 ( .A1(n2288), .A2(n2362), .ZN(n2398) );
  NAND2_X2 U88 ( .A1(n2286), .A2(n2642), .ZN(n2645) );
  NAND2_X2 U89 ( .A1(n2286), .A2(n2503), .ZN(n2506) );
  NAND2_X2 U90 ( .A1(n2286), .A2(n2362), .ZN(n2365) );
  NAND2_X2 U91 ( .A1(n2283), .A2(n2710), .ZN(n2712) );
  NAND2_X2 U92 ( .A1(n2283), .A2(n2605), .ZN(n2607) );
  NAND2_X2 U93 ( .A1(n2283), .A2(n2464), .ZN(n2466) );
  NAND2_X2 U94 ( .A1(n2283), .A2(n2323), .ZN(n2325) );
  NAND2_X2 U95 ( .A1(n2322), .A2(n2710), .ZN(n2678) );
  NAND2_X2 U96 ( .A1(n2322), .A2(n2605), .ZN(n2573) );
  NAND2_X2 U97 ( .A1(n2322), .A2(n2464), .ZN(n2432) );
  NAND2_X2 U98 ( .A1(n2284), .A2(n2283), .ZN(n2251) );
  AND2_X2 U99 ( .A1(n1648), .A2(n1652), .ZN(n1108) );
  AND2_X2 U100 ( .A1(n2238), .A2(n2243), .ZN(n1699) );
  AND2_X2 U101 ( .A1(n2236), .A2(n2243), .ZN(n1704) );
  AND2_X2 U102 ( .A1(n1646), .A2(n1652), .ZN(n1113) );
  AND2_X2 U103 ( .A1(n1648), .A2(n1653), .ZN(n1109) );
  AND2_X2 U104 ( .A1(n2238), .A2(n2242), .ZN(n1698) );
  AND2_X2 U105 ( .A1(n2236), .A2(n2242), .ZN(n1703) );
  AND2_X2 U106 ( .A1(n1646), .A2(n1653), .ZN(n1114) );
  AND2_X2 U107 ( .A1(n2227), .A2(n2242), .ZN(n1688) );
  AND2_X2 U108 ( .A1(n1637), .A2(n1652), .ZN(n1098) );
  NAND2_X2 U109 ( .A1(n1638), .A2(n1646), .ZN(n1089) );
  NAND2_X2 U110 ( .A1(n1638), .A2(n1643), .ZN(n1084) );
  NAND2_X2 U111 ( .A1(n1638), .A2(n1640), .ZN(n1079) );
  NAND2_X2 U112 ( .A1(n2228), .A2(n2236), .ZN(n1679) );
  NAND2_X2 U113 ( .A1(n2228), .A2(n2233), .ZN(n1674) );
  NAND2_X2 U114 ( .A1(n2228), .A2(n2230), .ZN(n1669) );
  NAND2_X2 U115 ( .A1(n1638), .A2(n1649), .ZN(n1094) );
  NAND2_X2 U116 ( .A1(n2228), .A2(n2239), .ZN(n1684) );
  NAND2_X2 U117 ( .A1(n2233), .A2(n2243), .ZN(n1694) );
  NAND2_X2 U118 ( .A1(n1643), .A2(n1653), .ZN(n1104) );
  NAND2_X2 U119 ( .A1(n2235), .A2(n2243), .ZN(n1706) );
  NAND2_X2 U120 ( .A1(n2230), .A2(n2243), .ZN(n1691) );
  NAND2_X2 U121 ( .A1(n2239), .A2(n2243), .ZN(n1701) );
  NAND2_X2 U122 ( .A1(n1645), .A2(n1653), .ZN(n1116) );
  NAND2_X2 U123 ( .A1(n1649), .A2(n1653), .ZN(n1111) );
  NAND2_X2 U124 ( .A1(n1640), .A2(n1653), .ZN(n1101) );
  NAND2_X2 U125 ( .A1(n2229), .A2(n2239), .ZN(n1683) );
  NAND2_X2 U126 ( .A1(n2229), .A2(n2233), .ZN(n1673) );
  NAND2_X2 U127 ( .A1(n2229), .A2(n2230), .ZN(n1668) );
  NAND2_X2 U128 ( .A1(n2229), .A2(n2236), .ZN(n1678) );
  NAND2_X2 U129 ( .A1(n1639), .A2(n1649), .ZN(n1093) );
  NAND2_X2 U130 ( .A1(n1639), .A2(n1646), .ZN(n1088) );
  NAND2_X2 U131 ( .A1(n1639), .A2(n1643), .ZN(n1083) );
  NAND2_X2 U132 ( .A1(n1639), .A2(n1640), .ZN(n1078) );
  NAND2_X2 U133 ( .A1(n1643), .A2(n1652), .ZN(n1103) );
  NAND2_X2 U134 ( .A1(n2233), .A2(n2242), .ZN(n1693) );
  NAND2_X2 U135 ( .A1(n1645), .A2(n1652), .ZN(n1117) );
  NAND2_X2 U136 ( .A1(n1649), .A2(n1652), .ZN(n1112) );
  NAND2_X2 U137 ( .A1(n1640), .A2(n1652), .ZN(n1102) );
  NAND2_X2 U138 ( .A1(n2235), .A2(n2242), .ZN(n1707) );
  NAND2_X2 U139 ( .A1(n2239), .A2(n2242), .ZN(n1702) );
  NAND2_X2 U140 ( .A1(n2230), .A2(n2242), .ZN(n1692) );
  AND2_X2 U141 ( .A1(n1639), .A2(n1637), .ZN(n1081) );
  AND2_X2 U142 ( .A1(n1639), .A2(n1648), .ZN(n1096) );
  AND2_X2 U143 ( .A1(n1639), .A2(n1645), .ZN(n1091) );
  AND2_X2 U144 ( .A1(n1639), .A2(n1642), .ZN(n1086) );
  AND2_X2 U145 ( .A1(n2228), .A2(n2227), .ZN(n1672) );
  AND2_X2 U146 ( .A1(n2238), .A2(n2228), .ZN(n1687) );
  AND2_X2 U147 ( .A1(n2228), .A2(n2235), .ZN(n1682) );
  AND2_X2 U148 ( .A1(n2228), .A2(n2232), .ZN(n1677) );
  AND2_X2 U149 ( .A1(n1642), .A2(n1652), .ZN(n1106) );
  AND2_X2 U150 ( .A1(n2232), .A2(n2243), .ZN(n1697) );
  AND2_X2 U151 ( .A1(n1638), .A2(n1637), .ZN(n1082) );
  AND2_X2 U152 ( .A1(n1648), .A2(n1638), .ZN(n1097) );
  AND2_X2 U153 ( .A1(n1638), .A2(n1645), .ZN(n1092) );
  AND2_X2 U154 ( .A1(n1638), .A2(n1642), .ZN(n1087) );
  AND2_X2 U155 ( .A1(n2229), .A2(n2238), .ZN(n1686) );
  AND2_X2 U156 ( .A1(n2229), .A2(n2227), .ZN(n1671) );
  AND2_X2 U157 ( .A1(n2229), .A2(n2235), .ZN(n1681) );
  AND2_X2 U158 ( .A1(n2229), .A2(n2232), .ZN(n1676) );
  AND2_X2 U159 ( .A1(n1642), .A2(n1653), .ZN(n1107) );
  AND2_X2 U160 ( .A1(n2232), .A2(n2242), .ZN(n1696) );
endmodule


module ImmGen ( instr, imm_out );
  input [31:0] instr;
  output [31:0] imm_out;
  wire   n24, n25, n26, n27, n28, n29, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n47;

  NAND3_X1 U50 ( .A1(instr[12]), .A2(n43), .A3(instr[14]), .ZN(n29) );
  NAND2_X1 U2 ( .A1(n27), .A2(n28), .ZN(n25) );
  NAND2_X1 U3 ( .A1(n45), .A2(n29), .ZN(n24) );
  INV_X1 U4 ( .A(n25), .ZN(n45) );
  OAI22_X1 U5 ( .A1(n16), .A2(n43), .B1(n25), .B2(n35), .ZN(imm_out[1]) );
  OAI22_X1 U6 ( .A1(n14), .A2(n36), .B1(n24), .B2(n20), .ZN(imm_out[8]) );
  OAI22_X1 U7 ( .A1(n15), .A2(n35), .B1(n24), .B2(n19), .ZN(imm_out[9]) );
  OAI22_X1 U8 ( .A1(n14), .A2(n34), .B1(n24), .B2(n18), .ZN(imm_out[10]) );
  INV_X1 U9 ( .A(n26), .ZN(imm_out[21]) );
  OAI21_X1 U10 ( .B1(n16), .B2(n33), .A(n26), .ZN(imm_out[11]) );
  OAI21_X1 U11 ( .B1(n14), .B2(n32), .A(n26), .ZN(imm_out[12]) );
  OAI21_X1 U12 ( .B1(n14), .B2(n31), .A(n26), .ZN(imm_out[13]) );
  OAI21_X1 U13 ( .B1(n15), .B2(n22), .A(n26), .ZN(imm_out[14]) );
  OAI21_X1 U14 ( .B1(n16), .B2(n21), .A(n26), .ZN(imm_out[15]) );
  OAI21_X1 U15 ( .B1(n15), .B2(n20), .A(n26), .ZN(imm_out[16]) );
  OAI21_X1 U16 ( .B1(n19), .B2(n16), .A(n26), .ZN(imm_out[17]) );
  OAI21_X1 U17 ( .B1(n14), .B2(n18), .A(n26), .ZN(imm_out[18]) );
  NAND4_X1 U18 ( .A1(instr[31]), .A2(n27), .A3(n28), .A4(n29), .ZN(n26) );
  NOR2_X1 U19 ( .A1(instr[2]), .A2(instr[5]), .ZN(n27) );
  OAI22_X1 U20 ( .A1(n44), .A2(n14), .B1(n25), .B2(n36), .ZN(imm_out[0]) );
  INV_X1 U21 ( .A(instr[12]), .ZN(n44) );
  OAI22_X1 U22 ( .A1(n42), .A2(n15), .B1(n25), .B2(n34), .ZN(imm_out[2]) );
  INV_X1 U23 ( .A(instr[14]), .ZN(n42) );
  OAI22_X1 U24 ( .A1(n14), .A2(n41), .B1(n25), .B2(n33), .ZN(imm_out[3]) );
  INV_X1 U25 ( .A(instr[15]), .ZN(n41) );
  OAI22_X1 U26 ( .A1(n15), .A2(n40), .B1(n25), .B2(n32), .ZN(imm_out[4]) );
  INV_X1 U27 ( .A(instr[16]), .ZN(n40) );
  OAI22_X1 U28 ( .A1(n15), .A2(n39), .B1(n25), .B2(n31), .ZN(imm_out[5]) );
  INV_X1 U29 ( .A(instr[17]), .ZN(n39) );
  OAI22_X1 U30 ( .A1(n16), .A2(n38), .B1(n24), .B2(n22), .ZN(imm_out[6]) );
  INV_X1 U31 ( .A(instr[18]), .ZN(n38) );
  OAI22_X1 U32 ( .A1(n16), .A2(n37), .B1(n24), .B2(n21), .ZN(imm_out[7]) );
  INV_X1 U33 ( .A(instr[19]), .ZN(n37) );
  OAI21_X1 U39 ( .B1(n15), .B2(n17), .A(n26), .ZN(imm_out[19]) );
  INV_X1 U40 ( .A(instr[31]), .ZN(n17) );
  INV_X1 U41 ( .A(instr[13]), .ZN(n43) );
  INV_X1 U42 ( .A(instr[21]), .ZN(n35) );
  INV_X1 U43 ( .A(instr[22]), .ZN(n34) );
  INV_X1 U44 ( .A(instr[23]), .ZN(n33) );
  INV_X1 U45 ( .A(instr[24]), .ZN(n32) );
  INV_X1 U46 ( .A(instr[20]), .ZN(n36) );
  INV_X1 U47 ( .A(instr[30]), .ZN(n18) );
  INV_X1 U48 ( .A(instr[25]), .ZN(n31) );
  INV_X1 U49 ( .A(instr[26]), .ZN(n22) );
  INV_X1 U52 ( .A(instr[27]), .ZN(n21) );
  INV_X1 U53 ( .A(instr[28]), .ZN(n20) );
  INV_X1 U54 ( .A(instr[29]), .ZN(n19) );
  INV_X1 U55 ( .A(n26), .ZN(imm_out[22]) );
  INV_X1 U56 ( .A(n26), .ZN(imm_out[23]) );
  INV_X1 U57 ( .A(n26), .ZN(imm_out[24]) );
  INV_X1 U58 ( .A(n26), .ZN(imm_out[25]) );
  INV_X1 U59 ( .A(n26), .ZN(imm_out[26]) );
  INV_X1 U60 ( .A(n26), .ZN(imm_out[27]) );
  INV_X1 U61 ( .A(n26), .ZN(imm_out[28]) );
  INV_X1 U62 ( .A(n26), .ZN(imm_out[29]) );
  INV_X1 U63 ( .A(n26), .ZN(imm_out[30]) );
  INV_X1 U64 ( .A(n26), .ZN(imm_out[31]) );
  INV_X1 U65 ( .A(n26), .ZN(imm_out[20]) );
  NAND3_X1 U34 ( .A1(n28), .A2(instr[5]), .A3(instr[2]), .ZN(n15) );
  NAND3_X1 U35 ( .A1(n28), .A2(instr[5]), .A3(instr[2]), .ZN(n14) );
  NAND3_X1 U36 ( .A1(n28), .A2(instr[5]), .A3(instr[2]), .ZN(n16) );
  NOR3_X1 U37 ( .A1(instr[6]), .A2(instr[3]), .A3(n47), .ZN(n28) );
  NAND3_X1 U38 ( .A1(instr[0]), .A2(instr[1]), .A3(instr[4]), .ZN(n47) );
endmodule


module control ( opcode, ALUsrc, ALUOP, regwrite, memtoreg, memread, memwrite, 
        branch );
  input [6:0] opcode;
  output [1:0] ALUOP;
  output ALUsrc, regwrite, memtoreg, memread, memwrite, branch;
  wire   n3, n4, n6, n14, n15;

  NAND4_X1 U9 ( .A1(opcode[4]), .A2(opcode[1]), .A3(n6), .A4(opcode[0]), .ZN(
        n4) );
  NOR2_X1 U12 ( .A1(opcode[6]), .A2(opcode[3]), .ZN(n6) );
  NOR2_X1 U13 ( .A1(n4), .A2(opcode[2]), .ZN(ALUOP[1]) );
  INV_X1 U15 ( .A(n3), .ZN(regwrite) );
  AOI21_X1 U16 ( .B1(n14), .B2(opcode[5]), .A(ALUOP[1]), .ZN(n3) );
  CLKBUF_X1 U17 ( .A(ALUsrc), .Z(ALUOP[0]) );
  INV_X1 U11 ( .A(n4), .ZN(n14) );
  NOR2_X1 U14 ( .A1(n4), .A2(n15), .ZN(ALUsrc) );
  XOR2_X1 U18 ( .A(opcode[2]), .B(opcode[5]), .Z(n15) );
endmodule


module REG_EX ( clk, rda, rdb, imm, wa, funct7, funct3, ALUsrc, ALUOP, 
        regwrite, branch, memread, memwrite, memtoreg, ra1, ra2, rda_EX, 
        rdb_EX, imm_EX, wa_EX, funct7_EX, funct3_EX, ALUsrc_EX, ALUOP_EX, 
        regwrite_EX, branch_EX, memread_EX, memwrite_EX, memtoreg_EX, ra1_EX, 
        ra2_EX );
  input [31:0] rda;
  input [31:0] rdb;
  input [31:0] imm;
  input [4:0] wa;
  input [2:0] funct3;
  input [1:0] ALUOP;
  input [4:0] ra1;
  input [4:0] ra2;
  output [31:0] rda_EX;
  output [31:0] rdb_EX;
  output [31:0] imm_EX;
  output [4:0] wa_EX;
  output [2:0] funct3_EX;
  output [1:0] ALUOP_EX;
  output [4:0] ra1_EX;
  output [4:0] ra2_EX;
  input clk, funct7, ALUsrc, regwrite, branch, memread, memwrite, memtoreg;
  output funct7_EX, ALUsrc_EX, regwrite_EX, branch_EX, memread_EX, memwrite_EX,
         memtoreg_EX;


  DFF_X1 rda_EX_reg_31_ ( .D(rda[31]), .CK(clk), .Q(rda_EX[31]) );
  DFF_X1 rda_EX_reg_30_ ( .D(rda[30]), .CK(clk), .Q(rda_EX[30]) );
  DFF_X1 rda_EX_reg_29_ ( .D(rda[29]), .CK(clk), .Q(rda_EX[29]) );
  DFF_X1 rda_EX_reg_28_ ( .D(rda[28]), .CK(clk), .Q(rda_EX[28]) );
  DFF_X1 rda_EX_reg_27_ ( .D(rda[27]), .CK(clk), .Q(rda_EX[27]) );
  DFF_X1 rda_EX_reg_26_ ( .D(rda[26]), .CK(clk), .Q(rda_EX[26]) );
  DFF_X1 rda_EX_reg_25_ ( .D(rda[25]), .CK(clk), .Q(rda_EX[25]) );
  DFF_X1 rda_EX_reg_24_ ( .D(rda[24]), .CK(clk), .Q(rda_EX[24]) );
  DFF_X1 rda_EX_reg_23_ ( .D(rda[23]), .CK(clk), .Q(rda_EX[23]) );
  DFF_X1 rda_EX_reg_22_ ( .D(rda[22]), .CK(clk), .Q(rda_EX[22]) );
  DFF_X1 rda_EX_reg_21_ ( .D(rda[21]), .CK(clk), .Q(rda_EX[21]) );
  DFF_X1 rda_EX_reg_20_ ( .D(rda[20]), .CK(clk), .Q(rda_EX[20]) );
  DFF_X1 rda_EX_reg_19_ ( .D(rda[19]), .CK(clk), .Q(rda_EX[19]) );
  DFF_X1 rda_EX_reg_18_ ( .D(rda[18]), .CK(clk), .Q(rda_EX[18]) );
  DFF_X1 rda_EX_reg_17_ ( .D(rda[17]), .CK(clk), .Q(rda_EX[17]) );
  DFF_X1 rda_EX_reg_16_ ( .D(rda[16]), .CK(clk), .Q(rda_EX[16]) );
  DFF_X1 rda_EX_reg_15_ ( .D(rda[15]), .CK(clk), .Q(rda_EX[15]) );
  DFF_X1 rda_EX_reg_14_ ( .D(rda[14]), .CK(clk), .Q(rda_EX[14]) );
  DFF_X1 rda_EX_reg_13_ ( .D(rda[13]), .CK(clk), .Q(rda_EX[13]) );
  DFF_X1 rda_EX_reg_12_ ( .D(rda[12]), .CK(clk), .Q(rda_EX[12]) );
  DFF_X1 rda_EX_reg_11_ ( .D(rda[11]), .CK(clk), .Q(rda_EX[11]) );
  DFF_X1 rda_EX_reg_10_ ( .D(rda[10]), .CK(clk), .Q(rda_EX[10]) );
  DFF_X1 rda_EX_reg_9_ ( .D(rda[9]), .CK(clk), .Q(rda_EX[9]) );
  DFF_X1 rda_EX_reg_8_ ( .D(rda[8]), .CK(clk), .Q(rda_EX[8]) );
  DFF_X1 rda_EX_reg_7_ ( .D(rda[7]), .CK(clk), .Q(rda_EX[7]) );
  DFF_X1 rda_EX_reg_6_ ( .D(rda[6]), .CK(clk), .Q(rda_EX[6]) );
  DFF_X1 rda_EX_reg_5_ ( .D(rda[5]), .CK(clk), .Q(rda_EX[5]) );
  DFF_X1 rda_EX_reg_4_ ( .D(rda[4]), .CK(clk), .Q(rda_EX[4]) );
  DFF_X1 rda_EX_reg_3_ ( .D(rda[3]), .CK(clk), .Q(rda_EX[3]) );
  DFF_X1 rda_EX_reg_2_ ( .D(rda[2]), .CK(clk), .Q(rda_EX[2]) );
  DFF_X1 rda_EX_reg_1_ ( .D(rda[1]), .CK(clk), .Q(rda_EX[1]) );
  DFF_X1 rda_EX_reg_0_ ( .D(rda[0]), .CK(clk), .Q(rda_EX[0]) );
  DFF_X1 rdb_EX_reg_31_ ( .D(rdb[31]), .CK(clk), .Q(rdb_EX[31]) );
  DFF_X1 rdb_EX_reg_30_ ( .D(rdb[30]), .CK(clk), .Q(rdb_EX[30]) );
  DFF_X1 rdb_EX_reg_29_ ( .D(rdb[29]), .CK(clk), .Q(rdb_EX[29]) );
  DFF_X1 rdb_EX_reg_28_ ( .D(rdb[28]), .CK(clk), .Q(rdb_EX[28]) );
  DFF_X1 rdb_EX_reg_27_ ( .D(rdb[27]), .CK(clk), .Q(rdb_EX[27]) );
  DFF_X1 rdb_EX_reg_26_ ( .D(rdb[26]), .CK(clk), .Q(rdb_EX[26]) );
  DFF_X1 rdb_EX_reg_25_ ( .D(rdb[25]), .CK(clk), .Q(rdb_EX[25]) );
  DFF_X1 rdb_EX_reg_24_ ( .D(rdb[24]), .CK(clk), .Q(rdb_EX[24]) );
  DFF_X1 rdb_EX_reg_23_ ( .D(rdb[23]), .CK(clk), .Q(rdb_EX[23]) );
  DFF_X1 rdb_EX_reg_22_ ( .D(rdb[22]), .CK(clk), .Q(rdb_EX[22]) );
  DFF_X1 rdb_EX_reg_21_ ( .D(rdb[21]), .CK(clk), .Q(rdb_EX[21]) );
  DFF_X1 rdb_EX_reg_20_ ( .D(rdb[20]), .CK(clk), .Q(rdb_EX[20]) );
  DFF_X1 rdb_EX_reg_19_ ( .D(rdb[19]), .CK(clk), .Q(rdb_EX[19]) );
  DFF_X1 rdb_EX_reg_18_ ( .D(rdb[18]), .CK(clk), .Q(rdb_EX[18]) );
  DFF_X1 rdb_EX_reg_17_ ( .D(rdb[17]), .CK(clk), .Q(rdb_EX[17]) );
  DFF_X1 rdb_EX_reg_16_ ( .D(rdb[16]), .CK(clk), .Q(rdb_EX[16]) );
  DFF_X1 rdb_EX_reg_15_ ( .D(rdb[15]), .CK(clk), .Q(rdb_EX[15]) );
  DFF_X1 rdb_EX_reg_14_ ( .D(rdb[14]), .CK(clk), .Q(rdb_EX[14]) );
  DFF_X1 rdb_EX_reg_13_ ( .D(rdb[13]), .CK(clk), .Q(rdb_EX[13]) );
  DFF_X1 rdb_EX_reg_12_ ( .D(rdb[12]), .CK(clk), .Q(rdb_EX[12]) );
  DFF_X1 rdb_EX_reg_11_ ( .D(rdb[11]), .CK(clk), .Q(rdb_EX[11]) );
  DFF_X1 rdb_EX_reg_10_ ( .D(rdb[10]), .CK(clk), .Q(rdb_EX[10]) );
  DFF_X1 rdb_EX_reg_9_ ( .D(rdb[9]), .CK(clk), .Q(rdb_EX[9]) );
  DFF_X1 rdb_EX_reg_8_ ( .D(rdb[8]), .CK(clk), .Q(rdb_EX[8]) );
  DFF_X1 rdb_EX_reg_7_ ( .D(rdb[7]), .CK(clk), .Q(rdb_EX[7]) );
  DFF_X1 rdb_EX_reg_6_ ( .D(rdb[6]), .CK(clk), .Q(rdb_EX[6]) );
  DFF_X1 rdb_EX_reg_5_ ( .D(rdb[5]), .CK(clk), .Q(rdb_EX[5]) );
  DFF_X1 rdb_EX_reg_4_ ( .D(rdb[4]), .CK(clk), .Q(rdb_EX[4]) );
  DFF_X1 rdb_EX_reg_3_ ( .D(rdb[3]), .CK(clk), .Q(rdb_EX[3]) );
  DFF_X1 rdb_EX_reg_2_ ( .D(rdb[2]), .CK(clk), .Q(rdb_EX[2]) );
  DFF_X1 rdb_EX_reg_1_ ( .D(rdb[1]), .CK(clk), .Q(rdb_EX[1]) );
  DFF_X1 rdb_EX_reg_0_ ( .D(rdb[0]), .CK(clk), .Q(rdb_EX[0]) );
  DFF_X1 imm_EX_reg_31_ ( .D(imm[31]), .CK(clk), .Q(imm_EX[31]) );
  DFF_X1 imm_EX_reg_30_ ( .D(imm[30]), .CK(clk), .Q(imm_EX[30]) );
  DFF_X1 imm_EX_reg_29_ ( .D(imm[29]), .CK(clk), .Q(imm_EX[29]) );
  DFF_X1 imm_EX_reg_28_ ( .D(imm[28]), .CK(clk), .Q(imm_EX[28]) );
  DFF_X1 imm_EX_reg_27_ ( .D(imm[27]), .CK(clk), .Q(imm_EX[27]) );
  DFF_X1 imm_EX_reg_26_ ( .D(imm[26]), .CK(clk), .Q(imm_EX[26]) );
  DFF_X1 imm_EX_reg_25_ ( .D(imm[25]), .CK(clk), .Q(imm_EX[25]) );
  DFF_X1 imm_EX_reg_24_ ( .D(imm[24]), .CK(clk), .Q(imm_EX[24]) );
  DFF_X1 imm_EX_reg_23_ ( .D(imm[23]), .CK(clk), .Q(imm_EX[23]) );
  DFF_X1 imm_EX_reg_22_ ( .D(imm[22]), .CK(clk), .Q(imm_EX[22]) );
  DFF_X1 imm_EX_reg_21_ ( .D(imm[21]), .CK(clk), .Q(imm_EX[21]) );
  DFF_X1 imm_EX_reg_20_ ( .D(imm[20]), .CK(clk), .Q(imm_EX[20]) );
  DFF_X1 imm_EX_reg_19_ ( .D(imm[19]), .CK(clk), .Q(imm_EX[19]) );
  DFF_X1 imm_EX_reg_18_ ( .D(imm[18]), .CK(clk), .Q(imm_EX[18]) );
  DFF_X1 imm_EX_reg_17_ ( .D(imm[17]), .CK(clk), .Q(imm_EX[17]) );
  DFF_X1 imm_EX_reg_16_ ( .D(imm[16]), .CK(clk), .Q(imm_EX[16]) );
  DFF_X1 imm_EX_reg_15_ ( .D(imm[15]), .CK(clk), .Q(imm_EX[15]) );
  DFF_X1 imm_EX_reg_14_ ( .D(imm[14]), .CK(clk), .Q(imm_EX[14]) );
  DFF_X1 imm_EX_reg_13_ ( .D(imm[13]), .CK(clk), .Q(imm_EX[13]) );
  DFF_X1 imm_EX_reg_12_ ( .D(imm[12]), .CK(clk), .Q(imm_EX[12]) );
  DFF_X1 imm_EX_reg_11_ ( .D(imm[11]), .CK(clk), .Q(imm_EX[11]) );
  DFF_X1 imm_EX_reg_10_ ( .D(imm[10]), .CK(clk), .Q(imm_EX[10]) );
  DFF_X1 imm_EX_reg_9_ ( .D(imm[9]), .CK(clk), .Q(imm_EX[9]) );
  DFF_X1 imm_EX_reg_8_ ( .D(imm[8]), .CK(clk), .Q(imm_EX[8]) );
  DFF_X1 imm_EX_reg_7_ ( .D(imm[7]), .CK(clk), .Q(imm_EX[7]) );
  DFF_X1 imm_EX_reg_6_ ( .D(imm[6]), .CK(clk), .Q(imm_EX[6]) );
  DFF_X1 imm_EX_reg_5_ ( .D(imm[5]), .CK(clk), .Q(imm_EX[5]) );
  DFF_X1 imm_EX_reg_4_ ( .D(imm[4]), .CK(clk), .Q(imm_EX[4]) );
  DFF_X1 imm_EX_reg_3_ ( .D(imm[3]), .CK(clk), .Q(imm_EX[3]) );
  DFF_X1 imm_EX_reg_2_ ( .D(imm[2]), .CK(clk), .Q(imm_EX[2]) );
  DFF_X1 imm_EX_reg_1_ ( .D(imm[1]), .CK(clk), .Q(imm_EX[1]) );
  DFF_X1 imm_EX_reg_0_ ( .D(imm[0]), .CK(clk), .Q(imm_EX[0]) );
  DFF_X1 wa_EX_reg_4_ ( .D(wa[4]), .CK(clk), .Q(wa_EX[4]) );
  DFF_X1 wa_EX_reg_3_ ( .D(wa[3]), .CK(clk), .Q(wa_EX[3]) );
  DFF_X1 wa_EX_reg_2_ ( .D(wa[2]), .CK(clk), .Q(wa_EX[2]) );
  DFF_X1 wa_EX_reg_1_ ( .D(wa[1]), .CK(clk), .Q(wa_EX[1]) );
  DFF_X1 wa_EX_reg_0_ ( .D(wa[0]), .CK(clk), .Q(wa_EX[0]) );
  DFF_X1 funct7_EX_reg ( .D(funct7), .CK(clk), .Q(funct7_EX) );
  DFF_X1 funct3_EX_reg_2_ ( .D(funct3[2]), .CK(clk), .Q(funct3_EX[2]) );
  DFF_X1 funct3_EX_reg_1_ ( .D(funct3[1]), .CK(clk), .Q(funct3_EX[1]) );
  DFF_X1 funct3_EX_reg_0_ ( .D(funct3[0]), .CK(clk), .Q(funct3_EX[0]) );
  DFF_X1 ALUsrc_EX_reg ( .D(ALUsrc), .CK(clk), .Q(ALUsrc_EX) );
  DFF_X1 ALUOP_EX_reg_1_ ( .D(ALUOP[1]), .CK(clk), .Q(ALUOP_EX[1]) );
  DFF_X1 ALUOP_EX_reg_0_ ( .D(ALUOP[0]), .CK(clk), .Q(ALUOP_EX[0]) );
  DFF_X1 regwrite_EX_reg ( .D(regwrite), .CK(clk), .Q(regwrite_EX) );
  DFF_X1 ra1_EX_reg_4_ ( .D(ra1[4]), .CK(clk), .Q(ra1_EX[4]) );
  DFF_X1 ra1_EX_reg_3_ ( .D(ra1[3]), .CK(clk), .Q(ra1_EX[3]) );
  DFF_X1 ra1_EX_reg_2_ ( .D(ra1[2]), .CK(clk), .Q(ra1_EX[2]) );
  DFF_X1 ra1_EX_reg_1_ ( .D(ra1[1]), .CK(clk), .Q(ra1_EX[1]) );
  DFF_X1 ra1_EX_reg_0_ ( .D(ra1[0]), .CK(clk), .Q(ra1_EX[0]) );
  DFF_X1 ra2_EX_reg_4_ ( .D(ra2[4]), .CK(clk), .Q(ra2_EX[4]) );
  DFF_X1 ra2_EX_reg_3_ ( .D(ra2[3]), .CK(clk), .Q(ra2_EX[3]) );
  DFF_X1 ra2_EX_reg_2_ ( .D(ra2[2]), .CK(clk), .Q(ra2_EX[2]) );
  DFF_X1 ra2_EX_reg_1_ ( .D(ra2[1]), .CK(clk), .Q(ra2_EX[1]) );
  DFF_X1 ra2_EX_reg_0_ ( .D(ra2[0]), .CK(clk), .Q(ra2_EX[0]) );
endmodule


module bit1adder_0 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n2;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n2), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n2) );
endmodule


module bit1adder_60 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_59 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N3 ( add1, add2, cin, result, cout );
  input [2:0] add1;
  input [2:0] add2;
  output [2:0] result;
  input cin;
  output cout;

  wire   [2:0] p;
  wire   [2:0] g;
  wire   [2:1] c_mid;

  XOR2_X1 U4 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U5 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U6 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_0 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), .sum(
        result[0]), .count(c_mid[1]) );
  bit1adder_60 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_59 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U2 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U3 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bit1adder_58 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_57 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_56 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_55 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N4_0 ( add1, add2, cin, result, cout );
  input [3:0] add1;
  input [3:0] add2;
  output [3:0] result;
  input cin;
  output cout;

  wire   [3:0] p;
  wire   [3:0] g;
  wire   [3:1] c_mid;

  XOR2_X1 U5 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U6 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U7 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U8 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_58 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), 
        .sum(result[0]), .count(c_mid[1]) );
  bit1adder_57 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_56 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_55 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U2 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U3 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U4 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bit1adder_54 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_53 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_52 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_51 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N4_1 ( add1, add2, cin, result, cout );
  input [3:0] add1;
  input [3:0] add2;
  output [3:0] result;
  input cin;
  output cout;

  wire   [3:0] p;
  wire   [3:0] g;
  wire   [3:1] c_mid;

  XOR2_X1 U5 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U6 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U7 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U8 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_54 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), 
        .sum(result[0]), .count(c_mid[1]) );
  bit1adder_53 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_52 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_51 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U2 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U3 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U4 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bitNmux_N4 ( in1, in0, sel, ou1 );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] ou1;
  input sel;
  wire   n7, n8, n9, n10, n11, n1;

  INV_X1 U1 ( .A(n11), .ZN(ou1[0]) );
  AOI22_X1 U2 ( .A1(in0[0]), .A2(n1), .B1(in1[0]), .B2(sel), .ZN(n11) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
  INV_X1 U4 ( .A(n8), .ZN(ou1[3]) );
  AOI22_X1 U5 ( .A1(in0[3]), .A2(n1), .B1(in1[3]), .B2(sel), .ZN(n8) );
  INV_X1 U6 ( .A(n7), .ZN(ou1[4]) );
  AOI22_X1 U7 ( .A1(in0[4]), .A2(n1), .B1(sel), .B2(in1[4]), .ZN(n7) );
  INV_X1 U8 ( .A(n9), .ZN(ou1[2]) );
  AOI22_X1 U9 ( .A1(in0[2]), .A2(n1), .B1(in1[2]), .B2(sel), .ZN(n9) );
  INV_X1 U10 ( .A(n10), .ZN(ou1[1]) );
  AOI22_X1 U11 ( .A1(in0[1]), .A2(n1), .B1(in1[1]), .B2(sel), .ZN(n10) );
endmodule


module bit1adder_50 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_49 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_48 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_47 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_46 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N5_0 ( add1, add2, cin, result, cout );
  input [4:0] add1;
  input [4:0] add2;
  output [4:0] result;
  input cin;
  output cout;

  wire   [4:0] p;
  wire   [4:0] g;
  wire   [4:1] c_mid;

  XOR2_X1 U6 ( .A(add2[4]), .B(add1[4]), .Z(p[4]) );
  XOR2_X1 U7 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U8 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U9 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U10 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_50 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), 
        .sum(result[0]), .count(c_mid[1]) );
  bit1adder_49 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_48 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_47 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(c_mid[4]) );
  bit1adder_46 block_4__bit1adder_module ( .g(g[4]), .p(p[4]), .cin(c_mid[4]), 
        .sum(result[4]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[4]), .A2(add1[4]), .ZN(g[4]) );
  AND2_X1 U2 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U3 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U4 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U5 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bit1adder_45 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_44 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_43 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_42 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_41 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N5_1 ( add1, add2, cin, result, cout );
  input [4:0] add1;
  input [4:0] add2;
  output [4:0] result;
  input cin;
  output cout;

  wire   [4:0] p;
  wire   [4:0] g;
  wire   [4:1] c_mid;

  XOR2_X1 U6 ( .A(add2[4]), .B(add1[4]), .Z(p[4]) );
  XOR2_X1 U7 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U8 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U9 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U10 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_45 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), 
        .sum(result[0]), .count(c_mid[1]) );
  bit1adder_44 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_43 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_42 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(c_mid[4]) );
  bit1adder_41 block_4__bit1adder_module ( .g(g[4]), .p(p[4]), .cin(c_mid[4]), 
        .sum(result[4]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[4]), .A2(add1[4]), .ZN(g[4]) );
  AND2_X1 U2 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U3 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U4 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U5 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bitNmux_N5 ( in1, in0, sel, ou1 );
  input [5:0] in1;
  input [5:0] in0;
  output [5:0] ou1;
  input sel;
  wire   n8, n9, n10, n11, n12, n13, n1;

  INV_X1 U1 ( .A(sel), .ZN(n1) );
  INV_X1 U2 ( .A(n13), .ZN(ou1[0]) );
  AOI22_X1 U3 ( .A1(in0[0]), .A2(n1), .B1(in1[0]), .B2(sel), .ZN(n13) );
  INV_X1 U4 ( .A(n8), .ZN(ou1[5]) );
  AOI22_X1 U5 ( .A1(in0[5]), .A2(n1), .B1(sel), .B2(in1[5]), .ZN(n8) );
  INV_X1 U6 ( .A(n10), .ZN(ou1[3]) );
  AOI22_X1 U7 ( .A1(in0[3]), .A2(n1), .B1(in1[3]), .B2(sel), .ZN(n10) );
  INV_X1 U8 ( .A(n9), .ZN(ou1[4]) );
  AOI22_X1 U9 ( .A1(in0[4]), .A2(n1), .B1(in1[4]), .B2(sel), .ZN(n9) );
  INV_X1 U10 ( .A(n11), .ZN(ou1[2]) );
  AOI22_X1 U11 ( .A1(in0[2]), .A2(n1), .B1(in1[2]), .B2(sel), .ZN(n11) );
  INV_X1 U12 ( .A(n12), .ZN(ou1[1]) );
  AOI22_X1 U13 ( .A1(in0[1]), .A2(n1), .B1(in1[1]), .B2(sel), .ZN(n12) );
endmodule


module bit1adder_40 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_39 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_38 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_37 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_36 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_35 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N6_0 ( add1, add2, cin, result, cout );
  input [5:0] add1;
  input [5:0] add2;
  output [5:0] result;
  input cin;
  output cout;

  wire   [5:0] p;
  wire   [5:0] g;
  wire   [5:1] c_mid;

  XOR2_X1 U7 ( .A(add2[5]), .B(add1[5]), .Z(p[5]) );
  XOR2_X1 U8 ( .A(add2[4]), .B(add1[4]), .Z(p[4]) );
  XOR2_X1 U9 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U10 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U11 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U12 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_40 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), 
        .sum(result[0]), .count(c_mid[1]) );
  bit1adder_39 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_38 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_37 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(c_mid[4]) );
  bit1adder_36 block_4__bit1adder_module ( .g(g[4]), .p(p[4]), .cin(c_mid[4]), 
        .sum(result[4]), .count(c_mid[5]) );
  bit1adder_35 block_5__bit1adder_module ( .g(g[5]), .p(p[5]), .cin(c_mid[5]), 
        .sum(result[5]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[5]), .A2(add1[5]), .ZN(g[5]) );
  AND2_X1 U2 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U3 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U4 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U5 ( .A1(add2[4]), .A2(add1[4]), .ZN(g[4]) );
  AND2_X1 U6 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bit1adder_34 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_33 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_32 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_31 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_30 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_29 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N6_1 ( add1, add2, cin, result, cout );
  input [5:0] add1;
  input [5:0] add2;
  output [5:0] result;
  input cin;
  output cout;

  wire   [5:0] p;
  wire   [5:0] g;
  wire   [5:1] c_mid;

  XOR2_X1 U7 ( .A(add2[5]), .B(add1[5]), .Z(p[5]) );
  XOR2_X1 U8 ( .A(add2[4]), .B(add1[4]), .Z(p[4]) );
  XOR2_X1 U9 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U10 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U11 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U12 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_34 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), 
        .sum(result[0]), .count(c_mid[1]) );
  bit1adder_33 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_32 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_31 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(c_mid[4]) );
  bit1adder_30 block_4__bit1adder_module ( .g(g[4]), .p(p[4]), .cin(c_mid[4]), 
        .sum(result[4]), .count(c_mid[5]) );
  bit1adder_29 block_5__bit1adder_module ( .g(g[5]), .p(p[5]), .cin(c_mid[5]), 
        .sum(result[5]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[5]), .A2(add1[5]), .ZN(g[5]) );
  AND2_X1 U2 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U3 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U4 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U5 ( .A1(add2[4]), .A2(add1[4]), .ZN(g[4]) );
  AND2_X1 U6 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bitNmux_N6 ( in1, in0, sel, ou1 );
  input [6:0] in1;
  input [6:0] in0;
  output [6:0] ou1;
  input sel;
  wire   n9, n10, n11, n12, n13, n14, n15, n1;

  INV_X1 U1 ( .A(sel), .ZN(n1) );
  INV_X1 U2 ( .A(n15), .ZN(ou1[0]) );
  AOI22_X1 U3 ( .A1(in0[0]), .A2(n1), .B1(in1[0]), .B2(sel), .ZN(n15) );
  INV_X1 U4 ( .A(n9), .ZN(ou1[6]) );
  AOI22_X1 U5 ( .A1(in0[6]), .A2(n1), .B1(sel), .B2(in1[6]), .ZN(n9) );
  INV_X1 U6 ( .A(n12), .ZN(ou1[3]) );
  AOI22_X1 U7 ( .A1(in0[3]), .A2(n1), .B1(in1[3]), .B2(sel), .ZN(n12) );
  INV_X1 U8 ( .A(n11), .ZN(ou1[4]) );
  AOI22_X1 U9 ( .A1(in0[4]), .A2(n1), .B1(in1[4]), .B2(sel), .ZN(n11) );
  INV_X1 U10 ( .A(n10), .ZN(ou1[5]) );
  AOI22_X1 U11 ( .A1(in0[5]), .A2(n1), .B1(in1[5]), .B2(sel), .ZN(n10) );
  INV_X1 U12 ( .A(n13), .ZN(ou1[2]) );
  AOI22_X1 U13 ( .A1(in0[2]), .A2(n1), .B1(in1[2]), .B2(sel), .ZN(n13) );
  INV_X1 U14 ( .A(n14), .ZN(ou1[1]) );
  AOI22_X1 U15 ( .A1(in0[1]), .A2(n1), .B1(in1[1]), .B2(sel), .ZN(n14) );
endmodule


module bit1adder_28 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_27 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_26 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_25 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_24 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_23 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_22 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N7_0 ( add1, add2, cin, result, cout );
  input [6:0] add1;
  input [6:0] add2;
  output [6:0] result;
  input cin;
  output cout;

  wire   [6:0] p;
  wire   [6:0] g;
  wire   [6:1] c_mid;

  XOR2_X1 U8 ( .A(add2[6]), .B(add1[6]), .Z(p[6]) );
  XOR2_X1 U9 ( .A(add2[5]), .B(add1[5]), .Z(p[5]) );
  XOR2_X1 U10 ( .A(add2[4]), .B(add1[4]), .Z(p[4]) );
  XOR2_X1 U11 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U12 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U13 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U14 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_28 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), 
        .sum(result[0]), .count(c_mid[1]) );
  bit1adder_27 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_26 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_25 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(c_mid[4]) );
  bit1adder_24 block_4__bit1adder_module ( .g(g[4]), .p(p[4]), .cin(c_mid[4]), 
        .sum(result[4]), .count(c_mid[5]) );
  bit1adder_23 block_5__bit1adder_module ( .g(g[5]), .p(p[5]), .cin(c_mid[5]), 
        .sum(result[5]), .count(c_mid[6]) );
  bit1adder_22 block_6__bit1adder_module ( .g(g[6]), .p(p[6]), .cin(c_mid[6]), 
        .sum(result[6]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[6]), .A2(add1[6]), .ZN(g[6]) );
  AND2_X1 U2 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U3 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U4 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U5 ( .A1(add2[4]), .A2(add1[4]), .ZN(g[4]) );
  AND2_X1 U6 ( .A1(add2[5]), .A2(add1[5]), .ZN(g[5]) );
  AND2_X1 U7 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bit1adder_21 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_20 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_19 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_18 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_17 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_16 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_15 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N7_3 ( add1, add2, cin, result, cout );
  input [6:0] add1;
  input [6:0] add2;
  output [6:0] result;
  input cin;
  output cout;

  wire   [6:0] p;
  wire   [6:0] g;
  wire   [6:1] c_mid;

  XOR2_X1 U8 ( .A(add2[6]), .B(add1[6]), .Z(p[6]) );
  XOR2_X1 U9 ( .A(add2[5]), .B(add1[5]), .Z(p[5]) );
  XOR2_X1 U10 ( .A(add2[4]), .B(add1[4]), .Z(p[4]) );
  XOR2_X1 U11 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U12 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U13 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U14 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_21 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), 
        .sum(result[0]), .count(c_mid[1]) );
  bit1adder_20 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_19 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_18 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(c_mid[4]) );
  bit1adder_17 block_4__bit1adder_module ( .g(g[4]), .p(p[4]), .cin(c_mid[4]), 
        .sum(result[4]), .count(c_mid[5]) );
  bit1adder_16 block_5__bit1adder_module ( .g(g[5]), .p(p[5]), .cin(c_mid[5]), 
        .sum(result[5]), .count(c_mid[6]) );
  bit1adder_15 block_6__bit1adder_module ( .g(g[6]), .p(p[6]), .cin(c_mid[6]), 
        .sum(result[6]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[6]), .A2(add1[6]), .ZN(g[6]) );
  AND2_X1 U2 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U3 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U4 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U5 ( .A1(add2[4]), .A2(add1[4]), .ZN(g[4]) );
  AND2_X1 U6 ( .A1(add2[5]), .A2(add1[5]), .ZN(g[5]) );
  AND2_X1 U7 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bitNmux_N7_0 ( in1, in0, sel, ou1 );
  input [7:0] in1;
  input [7:0] in0;
  output [7:0] ou1;
  input sel;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n1;

  INV_X1 U1 ( .A(sel), .ZN(n1) );
  INV_X1 U2 ( .A(n17), .ZN(ou1[0]) );
  AOI22_X1 U3 ( .A1(in0[0]), .A2(n1), .B1(in1[0]), .B2(sel), .ZN(n17) );
  INV_X1 U4 ( .A(n10), .ZN(ou1[7]) );
  AOI22_X1 U5 ( .A1(in0[7]), .A2(n1), .B1(sel), .B2(in1[7]), .ZN(n10) );
  INV_X1 U6 ( .A(n14), .ZN(ou1[3]) );
  AOI22_X1 U7 ( .A1(in0[3]), .A2(n1), .B1(in1[3]), .B2(sel), .ZN(n14) );
  INV_X1 U8 ( .A(n13), .ZN(ou1[4]) );
  AOI22_X1 U9 ( .A1(in0[4]), .A2(n1), .B1(in1[4]), .B2(sel), .ZN(n13) );
  INV_X1 U10 ( .A(n12), .ZN(ou1[5]) );
  AOI22_X1 U11 ( .A1(in0[5]), .A2(n1), .B1(in1[5]), .B2(sel), .ZN(n12) );
  INV_X1 U12 ( .A(n11), .ZN(ou1[6]) );
  AOI22_X1 U13 ( .A1(in0[6]), .A2(n1), .B1(in1[6]), .B2(sel), .ZN(n11) );
  INV_X1 U14 ( .A(n15), .ZN(ou1[2]) );
  AOI22_X1 U15 ( .A1(in0[2]), .A2(n1), .B1(in1[2]), .B2(sel), .ZN(n15) );
  INV_X1 U16 ( .A(n16), .ZN(ou1[1]) );
  AOI22_X1 U17 ( .A1(in0[1]), .A2(n1), .B1(in1[1]), .B2(sel), .ZN(n16) );
endmodule


module bit1adder_14 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_13 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_12 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_11 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_10 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_9 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_8 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N7_2 ( add1, add2, cin, result, cout );
  input [6:0] add1;
  input [6:0] add2;
  output [6:0] result;
  input cin;
  output cout;

  wire   [6:0] p;
  wire   [6:0] g;
  wire   [6:1] c_mid;

  XOR2_X1 U8 ( .A(add2[6]), .B(add1[6]), .Z(p[6]) );
  XOR2_X1 U9 ( .A(add2[5]), .B(add1[5]), .Z(p[5]) );
  XOR2_X1 U10 ( .A(add2[4]), .B(add1[4]), .Z(p[4]) );
  XOR2_X1 U11 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U12 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U13 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U14 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_14 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), 
        .sum(result[0]), .count(c_mid[1]) );
  bit1adder_13 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_12 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_11 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(c_mid[4]) );
  bit1adder_10 block_4__bit1adder_module ( .g(g[4]), .p(p[4]), .cin(c_mid[4]), 
        .sum(result[4]), .count(c_mid[5]) );
  bit1adder_9 block_5__bit1adder_module ( .g(g[5]), .p(p[5]), .cin(c_mid[5]), 
        .sum(result[5]), .count(c_mid[6]) );
  bit1adder_8 block_6__bit1adder_module ( .g(g[6]), .p(p[6]), .cin(c_mid[6]), 
        .sum(result[6]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[6]), .A2(add1[6]), .ZN(g[6]) );
  AND2_X1 U2 ( .A1(add2[5]), .A2(add1[5]), .ZN(g[5]) );
  AND2_X1 U3 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U4 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U5 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U6 ( .A1(add2[4]), .A2(add1[4]), .ZN(g[4]) );
  AND2_X1 U7 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bit1adder_7 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_6 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_5 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_4 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_3 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_2 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bit1adder_1 ( g, p, cin, sum, count );
  input g, p, cin;
  output sum, count;
  wire   n1;

  XOR2_X1 U3 ( .A(p), .B(cin), .Z(sum) );
  INV_X1 U1 ( .A(n1), .ZN(count) );
  AOI21_X1 U2 ( .B1(p), .B2(cin), .A(g), .ZN(n1) );
endmodule


module bitNRCAdder_N7_1 ( add1, add2, cin, result, cout );
  input [6:0] add1;
  input [6:0] add2;
  output [6:0] result;
  input cin;
  output cout;

  wire   [6:0] p;
  wire   [6:0] g;
  wire   [6:1] c_mid;

  XOR2_X1 U8 ( .A(add2[6]), .B(add1[6]), .Z(p[6]) );
  XOR2_X1 U9 ( .A(add2[5]), .B(add1[5]), .Z(p[5]) );
  XOR2_X1 U10 ( .A(add2[4]), .B(add1[4]), .Z(p[4]) );
  XOR2_X1 U11 ( .A(add2[3]), .B(add1[3]), .Z(p[3]) );
  XOR2_X1 U12 ( .A(add2[2]), .B(add1[2]), .Z(p[2]) );
  XOR2_X1 U13 ( .A(add2[1]), .B(add1[1]), .Z(p[1]) );
  XOR2_X1 U14 ( .A(add2[0]), .B(add1[0]), .Z(p[0]) );
  bit1adder_7 block_0__bit1adder_module ( .g(g[0]), .p(p[0]), .cin(cin), .sum(
        result[0]), .count(c_mid[1]) );
  bit1adder_6 block_1__bit1adder_module ( .g(g[1]), .p(p[1]), .cin(c_mid[1]), 
        .sum(result[1]), .count(c_mid[2]) );
  bit1adder_5 block_2__bit1adder_module ( .g(g[2]), .p(p[2]), .cin(c_mid[2]), 
        .sum(result[2]), .count(c_mid[3]) );
  bit1adder_4 block_3__bit1adder_module ( .g(g[3]), .p(p[3]), .cin(c_mid[3]), 
        .sum(result[3]), .count(c_mid[4]) );
  bit1adder_3 block_4__bit1adder_module ( .g(g[4]), .p(p[4]), .cin(c_mid[4]), 
        .sum(result[4]), .count(c_mid[5]) );
  bit1adder_2 block_5__bit1adder_module ( .g(g[5]), .p(p[5]), .cin(c_mid[5]), 
        .sum(result[5]), .count(c_mid[6]) );
  bit1adder_1 block_6__bit1adder_module ( .g(g[6]), .p(p[6]), .cin(c_mid[6]), 
        .sum(result[6]), .count(cout) );
  AND2_X1 U1 ( .A1(add2[6]), .A2(add1[6]), .ZN(g[6]) );
  AND2_X1 U2 ( .A1(add2[5]), .A2(add1[5]), .ZN(g[5]) );
  AND2_X1 U3 ( .A1(add2[1]), .A2(add1[1]), .ZN(g[1]) );
  AND2_X1 U4 ( .A1(add2[2]), .A2(add1[2]), .ZN(g[2]) );
  AND2_X1 U5 ( .A1(add2[3]), .A2(add1[3]), .ZN(g[3]) );
  AND2_X1 U6 ( .A1(add2[4]), .A2(add1[4]), .ZN(g[4]) );
  AND2_X1 U7 ( .A1(add2[0]), .A2(add1[0]), .ZN(g[0]) );
endmodule


module bitNmux_N7_1 ( in1, in0, sel, ou1 );
  input [7:0] in1;
  input [7:0] in0;
  output [7:0] ou1;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  INV_X1 U1 ( .A(sel), .ZN(n1) );
  AOI22_X1 U2 ( .A1(in0[0]), .A2(n1), .B1(in1[0]), .B2(sel), .ZN(n2) );
  INV_X1 U3 ( .A(n9), .ZN(ou1[7]) );
  AOI22_X1 U4 ( .A1(in0[7]), .A2(n1), .B1(sel), .B2(in1[7]), .ZN(n9) );
  INV_X1 U5 ( .A(n5), .ZN(ou1[3]) );
  AOI22_X1 U6 ( .A1(in0[3]), .A2(n1), .B1(in1[3]), .B2(sel), .ZN(n5) );
  INV_X1 U7 ( .A(n6), .ZN(ou1[4]) );
  AOI22_X1 U8 ( .A1(in0[4]), .A2(n1), .B1(in1[4]), .B2(sel), .ZN(n6) );
  INV_X1 U9 ( .A(n7), .ZN(ou1[5]) );
  AOI22_X1 U10 ( .A1(in0[5]), .A2(n1), .B1(in1[5]), .B2(sel), .ZN(n7) );
  INV_X1 U11 ( .A(n8), .ZN(ou1[6]) );
  AOI22_X1 U12 ( .A1(in0[6]), .A2(n1), .B1(in1[6]), .B2(sel), .ZN(n8) );
  INV_X1 U13 ( .A(n4), .ZN(ou1[2]) );
  AOI22_X1 U14 ( .A1(in0[2]), .A2(n1), .B1(in1[2]), .B2(sel), .ZN(n4) );
  INV_X1 U15 ( .A(n2), .ZN(ou1[0]) );
  INV_X1 U16 ( .A(n3), .ZN(ou1[1]) );
  AOI22_X1 U17 ( .A1(in0[1]), .A2(n1), .B1(in1[1]), .B2(sel), .ZN(n3) );
endmodule


module adder ( a, b, cin, sum, cout );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout;

  wire   [63:6] mid_sum;
  wire   [4:0] selected_c;
  wire   [9:0] mid_c;

  bitNRCAdder_N3 RCadder1_i1 ( .add1(a[2:0]), .add2(b[2:0]), .cin(cin), 
        .result(sum[2:0]), .cout(selected_c[0]) );
  bitNRCAdder_N4_0 RCadder1_i2 ( .add1(a[6:3]), .add2(b[6:3]), .cin(1'b0), 
        .result(mid_sum[9:6]), .cout(mid_c[0]) );
  bitNRCAdder_N4_1 RCadder2_i2 ( .add1(a[6:3]), .add2(b[6:3]), .cin(1'b1), 
        .result(mid_sum[13:10]), .cout(mid_c[1]) );
  bitNmux_N4 bit5mux_i2 ( .in1({mid_sum[13:10], mid_c[1]}), .in0({mid_sum[9:6], 
        mid_c[0]}), .sel(selected_c[0]), .ou1({sum[6:3], selected_c[1]}) );
  bitNRCAdder_N5_0 RCadder1_i3 ( .add1(a[11:7]), .add2(b[11:7]), .cin(1'b0), 
        .result(mid_sum[18:14]), .cout(mid_c[2]) );
  bitNRCAdder_N5_1 RCadder2_i3 ( .add1(a[11:7]), .add2(b[11:7]), .cin(1'b1), 
        .result(mid_sum[23:19]), .cout(mid_c[3]) );
  bitNmux_N5 bit5mux_i3 ( .in1({mid_sum[23:19], mid_c[3]}), .in0({
        mid_sum[18:14], mid_c[2]}), .sel(selected_c[1]), .ou1({sum[11:7], 
        selected_c[2]}) );
  bitNRCAdder_N6_0 RCadder1_i4 ( .add1(a[17:12]), .add2(b[17:12]), .cin(1'b0), 
        .result(mid_sum[29:24]), .cout(mid_c[4]) );
  bitNRCAdder_N6_1 RCadder2_i4 ( .add1(a[17:12]), .add2(b[17:12]), .cin(1'b1), 
        .result(mid_sum[35:30]), .cout(mid_c[5]) );
  bitNmux_N6 bit5mux_i4 ( .in1({mid_sum[35:30], mid_c[5]}), .in0({
        mid_sum[29:24], mid_c[4]}), .sel(selected_c[2]), .ou1({sum[17:12], 
        selected_c[3]}) );
  bitNRCAdder_N7_0 RCadder1_i5 ( .add1(a[24:18]), .add2(b[24:18]), .cin(1'b0), 
        .result(mid_sum[42:36]), .cout(mid_c[6]) );
  bitNRCAdder_N7_3 RCadder2_i5 ( .add1(a[24:18]), .add2(b[24:18]), .cin(1'b1), 
        .result(mid_sum[49:43]), .cout(mid_c[7]) );
  bitNmux_N7_0 bit5mux_i5 ( .in1({mid_sum[49:43], mid_c[7]}), .in0({
        mid_sum[42:36], mid_c[6]}), .sel(selected_c[3]), .ou1({sum[24:18], 
        selected_c[4]}) );
  bitNRCAdder_N7_2 RCadder1_i6 ( .add1(a[31:25]), .add2(b[31:25]), .cin(1'b0), 
        .result(mid_sum[56:50]), .cout(mid_c[8]) );
  bitNRCAdder_N7_1 RCadder2_i6 ( .add1(a[31:25]), .add2(b[31:25]), .cin(1'b1), 
        .result(mid_sum[63:57]), .cout(mid_c[9]) );
  bitNmux_N7_1 bit5mux_i6 ( .in1({mid_sum[63:57], mid_c[9]}), .in0({
        mid_sum[56:50], mid_c[8]}), .sel(selected_c[4]), .ou1({sum[31:25], 
        cout}) );
endmodule


module alu_32bit ( alu_src1, alu_src2, alu_control, alu_result );
  input [31:0] alu_src1;
  input [31:0] alu_src2;
  input [3:0] alu_control;
  output [31:0] alu_result;
  wire   adder_cout, sra_result_30_, sra_result_29_, sra_result_28_,
         sra_result_27_, sra_result_26_, sra_result_25_, sra_result_24_,
         sra_result_23_, sra_result_22_, sra_result_21_, sra_result_20_,
         sra_result_19_, sra_result_18_, sra_result_17_, sra_result_16_,
         sra_result_15_, sra_result_14_, sra_result_13_, sra_result_12_,
         sra_result_11_, sra_result_10_, sra_result_9_, sra_result_8_,
         sra_result_7_, sra_result_6_, sra_result_5_, sra_result_4_,
         sra_result_3_, sra_result_2_, sra_result_1_, sra_result_0_, N96, n46,
         n47, n48, n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n1, n2, n3, n4, n5, n6, n8, n11, n16, n17, n18, n22, n23,
         n25, n29, n31, n32, n33, n40, n41, n42, n43, n44, n45, n53, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n223, n224, n225, n226, n227, n229, n230,
         n231, n232, n235, n236, n237, n238, n239, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825;
  wire   [31:0] adder_operand2;
  wire   [31:0] adder_result;
  wire   [31:0] sll_result;
  wire   [31:0] srl_result;

  NAND3_X1 U214 ( .A1(n86), .A2(n87), .A3(n88), .ZN(alu_result[30]) );
  NAND3_X1 U215 ( .A1(n95), .A2(n96), .A3(n97), .ZN(alu_result[29]) );
  NAND3_X1 U216 ( .A1(n100), .A2(n101), .A3(n102), .ZN(alu_result[28]) );
  NAND3_X1 U217 ( .A1(n105), .A2(n106), .A3(n107), .ZN(alu_result[27]) );
  NAND3_X1 U218 ( .A1(n110), .A2(n111), .A3(n112), .ZN(alu_result[26]) );
  NAND3_X1 U219 ( .A1(n115), .A2(n116), .A3(n117), .ZN(alu_result[25]) );
  NAND3_X1 U220 ( .A1(n120), .A2(n121), .A3(n122), .ZN(alu_result[24]) );
  NAND3_X1 U221 ( .A1(n125), .A2(n126), .A3(n127), .ZN(alu_result[23]) );
  NAND3_X1 U222 ( .A1(n130), .A2(n131), .A3(n132), .ZN(alu_result[22]) );
  NAND3_X1 U223 ( .A1(n135), .A2(n136), .A3(n137), .ZN(alu_result[21]) );
  NAND3_X1 U224 ( .A1(n140), .A2(n141), .A3(n142), .ZN(alu_result[20]) );
  NAND3_X1 U225 ( .A1(n149), .A2(n150), .A3(n151), .ZN(alu_result[19]) );
  NAND3_X1 U226 ( .A1(n154), .A2(n155), .A3(n156), .ZN(alu_result[18]) );
  NAND3_X1 U227 ( .A1(n159), .A2(n160), .A3(n161), .ZN(alu_result[17]) );
  NAND3_X1 U228 ( .A1(n164), .A2(n165), .A3(n166), .ZN(alu_result[16]) );
  NAND3_X1 U229 ( .A1(n169), .A2(n170), .A3(n171), .ZN(alu_result[15]) );
  NAND3_X1 U230 ( .A1(n174), .A2(n175), .A3(n176), .ZN(alu_result[14]) );
  NAND3_X1 U231 ( .A1(n179), .A2(n180), .A3(n181), .ZN(alu_result[13]) );
  NAND3_X1 U232 ( .A1(n184), .A2(n185), .A3(n186), .ZN(alu_result[12]) );
  OAI33_X1 U233 ( .A1(n320), .A2(n53), .A3(n51), .B1(n201), .B2(n321), .B3(
        n322), .ZN(n200) );
  XOR2_X1 U236 ( .A(alu_src2[9]), .B(N96), .Z(adder_operand2[9]) );
  XOR2_X1 U237 ( .A(alu_src2[8]), .B(N96), .Z(adder_operand2[8]) );
  XOR2_X1 U238 ( .A(alu_src2[7]), .B(N96), .Z(adder_operand2[7]) );
  XOR2_X1 U239 ( .A(alu_src2[6]), .B(N96), .Z(adder_operand2[6]) );
  XOR2_X1 U240 ( .A(n239), .B(N96), .Z(adder_operand2[5]) );
  XOR2_X1 U241 ( .A(alu_src2[4]), .B(N96), .Z(adder_operand2[4]) );
  XOR2_X1 U242 ( .A(n216), .B(N96), .Z(adder_operand2[3]) );
  XOR2_X1 U243 ( .A(alu_src2[31]), .B(N96), .Z(adder_operand2[31]) );
  XOR2_X1 U244 ( .A(alu_src2[30]), .B(N96), .Z(adder_operand2[30]) );
  XOR2_X1 U245 ( .A(n211), .B(N96), .Z(adder_operand2[2]) );
  XOR2_X1 U246 ( .A(alu_src2[29]), .B(N96), .Z(adder_operand2[29]) );
  XOR2_X1 U247 ( .A(alu_src2[28]), .B(N96), .Z(adder_operand2[28]) );
  XOR2_X1 U248 ( .A(alu_src2[27]), .B(N96), .Z(adder_operand2[27]) );
  XOR2_X1 U249 ( .A(alu_src2[26]), .B(N96), .Z(adder_operand2[26]) );
  XOR2_X1 U250 ( .A(alu_src2[25]), .B(N96), .Z(adder_operand2[25]) );
  XOR2_X1 U251 ( .A(alu_src2[24]), .B(N96), .Z(adder_operand2[24]) );
  XOR2_X1 U252 ( .A(alu_src2[23]), .B(N96), .Z(adder_operand2[23]) );
  XOR2_X1 U253 ( .A(alu_src2[22]), .B(N96), .Z(adder_operand2[22]) );
  XOR2_X1 U254 ( .A(alu_src2[21]), .B(N96), .Z(adder_operand2[21]) );
  XOR2_X1 U255 ( .A(alu_src2[20]), .B(N96), .Z(adder_operand2[20]) );
  XOR2_X1 U256 ( .A(n206), .B(N96), .Z(adder_operand2[1]) );
  XOR2_X1 U257 ( .A(alu_src2[19]), .B(N96), .Z(adder_operand2[19]) );
  XOR2_X1 U258 ( .A(alu_src2[18]), .B(N96), .Z(adder_operand2[18]) );
  XOR2_X1 U259 ( .A(alu_src2[17]), .B(N96), .Z(adder_operand2[17]) );
  XOR2_X1 U260 ( .A(alu_src2[16]), .B(N96), .Z(adder_operand2[16]) );
  XOR2_X1 U261 ( .A(alu_src2[15]), .B(N96), .Z(adder_operand2[15]) );
  XOR2_X1 U262 ( .A(alu_src2[14]), .B(N96), .Z(adder_operand2[14]) );
  XOR2_X1 U263 ( .A(alu_src2[13]), .B(N96), .Z(adder_operand2[13]) );
  XOR2_X1 U264 ( .A(alu_src2[12]), .B(N96), .Z(adder_operand2[12]) );
  XOR2_X1 U265 ( .A(alu_src2[11]), .B(N96), .Z(adder_operand2[11]) );
  XOR2_X1 U266 ( .A(alu_src2[10]), .B(N96), .Z(adder_operand2[10]) );
  XOR2_X1 U267 ( .A(n44), .B(N96), .Z(adder_operand2[0]) );
  adder adder_module ( .a({n41, alu_src1[30:0]}), .b(adder_operand2), .cin(N96), .sum(adder_result), .cout(adder_cout) );
  CLKBUF_X1 U2 ( .A(n629), .Z(n11) );
  CLKBUF_X1 U3 ( .A(n476), .Z(n8) );
  CLKBUF_X1 U6 ( .A(alu_src2[5]), .Z(n238) );
  CLKBUF_X1 U7 ( .A(alu_src2[5]), .Z(n237) );
  CLKBUF_X1 U8 ( .A(alu_src2[5]), .Z(n235) );
  CLKBUF_X1 U9 ( .A(alu_src2[5]), .Z(n236) );
  NOR3_X1 U10 ( .A1(n434), .A2(n238), .A3(n8), .ZN(sll_result[27]) );
  INV_X1 U11 ( .A(n430), .ZN(n258) );
  NOR3_X1 U12 ( .A1(n624), .A2(n239), .A3(n11), .ZN(srl_result[8]) );
  NOR4_X1 U13 ( .A1(n237), .A2(alu_src2[4]), .A3(n629), .A4(n581), .ZN(
        srl_result[31]) );
  NOR4_X1 U14 ( .A1(n237), .A2(alu_src2[4]), .A3(n629), .A4(n567), .ZN(
        srl_result[27]) );
  NOR4_X1 U15 ( .A1(n237), .A2(alu_src2[4]), .A3(n629), .A4(n568), .ZN(
        srl_result[28]) );
  NOR4_X1 U16 ( .A1(n237), .A2(alu_src2[4]), .A3(n629), .A4(n569), .ZN(
        srl_result[29]) );
  NOR4_X1 U17 ( .A1(n237), .A2(alu_src2[4]), .A3(n629), .A4(n580), .ZN(
        srl_result[30]) );
  NOR4_X1 U18 ( .A1(n236), .A2(n225), .A3(n539), .A4(n629), .ZN(srl_result[16]) );
  NOR4_X1 U19 ( .A1(n236), .A2(n224), .A3(n553), .A4(n629), .ZN(srl_result[17]) );
  NOR4_X1 U20 ( .A1(n236), .A2(n224), .A3(n577), .A4(n11), .ZN(srl_result[18])
         );
  NOR4_X1 U21 ( .A1(n236), .A2(n224), .A3(n589), .A4(n629), .ZN(srl_result[19]) );
  NOR4_X1 U22 ( .A1(n236), .A2(n224), .A3(n596), .A4(n11), .ZN(srl_result[20])
         );
  NOR4_X1 U23 ( .A1(n236), .A2(n224), .A3(n603), .A4(n11), .ZN(srl_result[21])
         );
  NOR4_X1 U24 ( .A1(n236), .A2(n223), .A3(n610), .A4(n629), .ZN(srl_result[22]) );
  NOR4_X1 U25 ( .A1(n236), .A2(n223), .A3(n617), .A4(n11), .ZN(srl_result[23])
         );
  NOR4_X1 U26 ( .A1(n237), .A2(n223), .A3(n629), .A4(n622), .ZN(srl_result[24]) );
  NOR4_X1 U27 ( .A1(n237), .A2(n223), .A3(n629), .A4(n627), .ZN(srl_result[25]) );
  NOR4_X1 U28 ( .A1(n237), .A2(n223), .A3(n629), .A4(n566), .ZN(srl_result[26]) );
  NOR4_X1 U29 ( .A1(n235), .A2(n226), .A3(n476), .A4(n380), .ZN(sll_result[1])
         );
  NOR4_X1 U30 ( .A1(n236), .A2(n225), .A3(n476), .A4(n474), .ZN(sll_result[7])
         );
  NOR4_X1 U31 ( .A1(n236), .A2(n225), .A3(n475), .A4(n8), .ZN(sll_result[8])
         );
  NOR4_X1 U32 ( .A1(n236), .A2(n225), .A3(n477), .A4(n476), .ZN(sll_result[9])
         );
  NOR4_X1 U33 ( .A1(n235), .A2(n227), .A3(n432), .A4(n476), .ZN(sll_result[11]) );
  NOR4_X1 U34 ( .A1(n235), .A2(n227), .A3(n440), .A4(n8), .ZN(sll_result[12])
         );
  NOR4_X1 U35 ( .A1(n235), .A2(n227), .A3(n448), .A4(n8), .ZN(sll_result[13])
         );
  NOR4_X1 U36 ( .A1(n235), .A2(n227), .A3(n458), .A4(n476), .ZN(sll_result[14]) );
  NOR4_X1 U37 ( .A1(n235), .A2(n227), .A3(n467), .A4(n8), .ZN(sll_result[15])
         );
  NOR4_X1 U38 ( .A1(n235), .A2(alu_src2[4]), .A3(n476), .A4(n361), .ZN(
        sll_result[0]) );
  NOR4_X1 U39 ( .A1(n235), .A2(alu_src2[4]), .A3(n425), .A4(n476), .ZN(
        sll_result[10]) );
  NOR3_X1 U40 ( .A1(n363), .A2(n238), .A3(n476), .ZN(sll_result[16]) );
  NOR3_X1 U41 ( .A1(n379), .A2(n238), .A3(n8), .ZN(sll_result[19]) );
  NOR3_X1 U42 ( .A1(n392), .A2(n238), .A3(n8), .ZN(sll_result[21]) );
  NOR3_X1 U43 ( .A1(n398), .A2(n238), .A3(n8), .ZN(sll_result[22]) );
  NOR3_X1 U44 ( .A1(n404), .A2(n238), .A3(n8), .ZN(sll_result[23]) );
  NOR3_X1 U45 ( .A1(n427), .A2(n238), .A3(n8), .ZN(sll_result[26]) );
  INV_X1 U46 ( .A(n423), .ZN(n261) );
  INV_X1 U47 ( .A(n556), .ZN(n243) );
  INV_X1 U48 ( .A(n558), .ZN(n247) );
  INV_X1 U49 ( .A(n560), .ZN(n245) );
  INV_X1 U50 ( .A(n562), .ZN(n246) );
  INV_X1 U51 ( .A(n409), .ZN(n317) );
  INV_X1 U52 ( .A(n417), .ZN(n318) );
  INV_X1 U53 ( .A(n372), .ZN(n314) );
  INV_X1 U54 ( .A(n402), .ZN(n298) );
  NOR3_X1 U55 ( .A1(n630), .A2(n239), .A3(n11), .ZN(srl_result[9]) );
  NOR3_X1 U56 ( .A1(n507), .A2(n237), .A3(n11), .ZN(srl_result[10]) );
  NOR3_X1 U57 ( .A1(n513), .A2(n237), .A3(n11), .ZN(srl_result[11]) );
  NOR3_X1 U58 ( .A1(n518), .A2(n237), .A3(n11), .ZN(srl_result[12]) );
  NOR3_X1 U59 ( .A1(n526), .A2(n237), .A3(n11), .ZN(srl_result[13]) );
  NOR3_X1 U60 ( .A1(n531), .A2(n238), .A3(n11), .ZN(srl_result[14]) );
  NOR3_X1 U61 ( .A1(n538), .A2(n237), .A3(n11), .ZN(srl_result[15]) );
  NOR3_X1 U62 ( .A1(n450), .A2(n238), .A3(n8), .ZN(sll_result[29]) );
  INV_X1 U63 ( .A(n446), .ZN(n252) );
  NOR3_X1 U64 ( .A1(n368), .A2(n238), .A3(n8), .ZN(sll_result[17]) );
  NOR3_X1 U65 ( .A1(n374), .A2(n238), .A3(n8), .ZN(sll_result[18]) );
  NOR3_X1 U66 ( .A1(n386), .A2(n238), .A3(n8), .ZN(sll_result[20]) );
  NOR3_X1 U67 ( .A1(n442), .A2(n238), .A3(n8), .ZN(sll_result[28]) );
  INV_X1 U68 ( .A(n438), .ZN(n255) );
  OR2_X1 U69 ( .A1(n564), .A2(n217), .ZN(n622) );
  OR2_X1 U70 ( .A1(n565), .A2(n217), .ZN(n627) );
  OR2_X1 U71 ( .A1(n544), .A2(n216), .ZN(n566) );
  OR2_X1 U72 ( .A1(n546), .A2(n216), .ZN(n567) );
  OR2_X1 U73 ( .A1(n384), .A2(n218), .ZN(n471) );
  OR2_X1 U74 ( .A1(n390), .A2(alu_src2[3]), .ZN(n472) );
  OR2_X1 U75 ( .A1(n396), .A2(n217), .ZN(n473) );
  OR2_X1 U76 ( .A1(n524), .A2(n209), .ZN(n536) );
  INV_X1 U77 ( .A(n592), .ZN(n300) );
  INV_X1 U78 ( .A(n436), .ZN(n267) );
  INV_X1 U79 ( .A(n444), .ZN(n264) );
  INV_X1 U80 ( .A(n219), .ZN(n216) );
  INV_X1 U81 ( .A(n210), .ZN(n206) );
  INV_X1 U82 ( .A(n205), .ZN(n44) );
  CLKBUF_X2 U83 ( .A(alu_src2[5]), .Z(n239) );
  INV_X1 U84 ( .A(adder_result[31]), .ZN(n241) );
  INV_X1 U85 ( .A(n205), .ZN(n53) );
  INV_X1 U86 ( .A(n43), .ZN(n42) );
  NOR3_X1 U87 ( .A1(n629), .A2(n237), .A3(n492), .ZN(srl_result[0]) );
  INV_X1 U88 ( .A(n488), .ZN(n299) );
  INV_X1 U89 ( .A(n210), .ZN(n207) );
  INV_X1 U90 ( .A(n205), .ZN(n45) );
  NAND2_X1 U91 ( .A1(n145), .A2(n146), .ZN(alu_result[1]) );
  AOI222_X1 U92 ( .A1(adder_result[1]), .A2(n23), .B1(srl_result[1]), .B2(n54), 
        .C1(sll_result[1]), .C2(n17), .ZN(n145) );
  AOI221_X1 U93 ( .B1(sra_result_1_), .B2(n48), .C1(n206), .C2(n147), .A(n148), 
        .ZN(n146) );
  NAND2_X1 U94 ( .A1(n91), .A2(n92), .ZN(alu_result[2]) );
  AOI222_X1 U95 ( .A1(adder_result[2]), .A2(n22), .B1(srl_result[2]), .B2(n54), 
        .C1(sll_result[2]), .C2(n16), .ZN(n91) );
  AOI221_X1 U96 ( .B1(sra_result_2_), .B2(n48), .C1(n211), .C2(n93), .A(n94), 
        .ZN(n92) );
  NOR4_X1 U97 ( .A1(n235), .A2(n226), .A3(n476), .A4(n451), .ZN(sll_result[2])
         );
  NAND2_X1 U98 ( .A1(n72), .A2(n73), .ZN(alu_result[4]) );
  AOI222_X1 U99 ( .A1(adder_result[4]), .A2(n22), .B1(srl_result[4]), .B2(n54), 
        .C1(sll_result[4]), .C2(n16), .ZN(n72) );
  AOI221_X1 U100 ( .B1(sra_result_4_), .B2(n48), .C1(alu_src2[4]), .C2(n74), 
        .A(n75), .ZN(n73) );
  NOR4_X1 U101 ( .A1(n235), .A2(n226), .A3(n476), .A4(n471), .ZN(sll_result[4]) );
  NAND2_X1 U102 ( .A1(n68), .A2(n69), .ZN(alu_result[5]) );
  AOI222_X1 U103 ( .A1(adder_result[5]), .A2(n22), .B1(srl_result[5]), .B2(n54), .C1(sll_result[5]), .C2(n16), .ZN(n68) );
  AOI221_X1 U104 ( .B1(sra_result_5_), .B2(n48), .C1(n239), .C2(n70), .A(n71), 
        .ZN(n69) );
  NOR4_X1 U105 ( .A1(n235), .A2(n226), .A3(n476), .A4(n472), .ZN(sll_result[5]) );
  NOR3_X1 U106 ( .A1(n555), .A2(n238), .A3(n11), .ZN(srl_result[1]) );
  NAND2_X1 U107 ( .A1(n40), .A2(n205), .ZN(n524) );
  INV_X1 U108 ( .A(n500), .ZN(n271) );
  INV_X1 U109 ( .A(n490), .ZN(n244) );
  INV_X1 U110 ( .A(n339), .ZN(n288) );
  INV_X1 U111 ( .A(n210), .ZN(n208) );
  INV_X1 U112 ( .A(n43), .ZN(n40) );
  INV_X1 U113 ( .A(n43), .ZN(n41) );
  NOR3_X1 U114 ( .A1(n598), .A2(n239), .A3(n11), .ZN(srl_result[4]) );
  NOR3_X1 U115 ( .A1(n476), .A2(n238), .A3(n469), .ZN(sll_result[31]) );
  INV_X1 U116 ( .A(n465), .ZN(n242) );
  NOR3_X1 U117 ( .A1(n412), .A2(n238), .A3(n8), .ZN(sll_result[24]) );
  NOR3_X1 U118 ( .A1(n460), .A2(n238), .A3(n476), .ZN(sll_result[30]) );
  INV_X1 U119 ( .A(n456), .ZN(n249) );
  INV_X1 U120 ( .A(n210), .ZN(n209) );
  INV_X1 U121 ( .A(n219), .ZN(n217) );
  INV_X1 U122 ( .A(n219), .ZN(n218) );
  INV_X1 U123 ( .A(n205), .ZN(n204) );
  NOR2_X1 U124 ( .A1(n244), .A2(n211), .ZN(n556) );
  NOR2_X1 U125 ( .A1(n529), .A2(n211), .ZN(n560) );
  NOR2_X1 U126 ( .A1(n366), .A2(n211), .ZN(n417) );
  NOR2_X1 U127 ( .A1(n542), .A2(n211), .ZN(n558) );
  NOR2_X1 U128 ( .A1(n536), .A2(n211), .ZN(n562) );
  NOR2_X1 U129 ( .A1(n341), .A2(n211), .ZN(n409) );
  NOR2_X1 U130 ( .A1(n351), .A2(n211), .ZN(n372) );
  CLKBUF_X1 U131 ( .A(alu_src2[4]), .Z(n229) );
  CLKBUF_X1 U132 ( .A(alu_src2[4]), .Z(n230) );
  CLKBUF_X1 U133 ( .A(alu_src2[4]), .Z(n231) );
  CLKBUF_X1 U135 ( .A(alu_src2[4]), .Z(n232) );
  NAND2_X1 U140 ( .A1(n556), .A2(n219), .ZN(n568) );
  NAND2_X1 U141 ( .A1(n558), .A2(n219), .ZN(n569) );
  NAND2_X1 U142 ( .A1(n560), .A2(n219), .ZN(n580) );
  NAND2_X1 U143 ( .A1(n562), .A2(n219), .ZN(n581) );
  NAND2_X1 U144 ( .A1(n409), .A2(n219), .ZN(n361) );
  NAND2_X1 U145 ( .A1(n417), .A2(n219), .ZN(n380) );
  NAND2_X1 U146 ( .A1(n372), .A2(n219), .ZN(n451) );
  NAND2_X1 U147 ( .A1(n402), .A2(n219), .ZN(n474) );
  NOR3_X1 U150 ( .A1(n579), .A2(n238), .A3(n11), .ZN(srl_result[2]) );
  NOR3_X1 U151 ( .A1(n591), .A2(n238), .A3(n11), .ZN(srl_result[3]) );
  NOR3_X1 U152 ( .A1(n605), .A2(n238), .A3(n11), .ZN(srl_result[5]) );
  NOR3_X1 U153 ( .A1(n612), .A2(n239), .A3(n629), .ZN(srl_result[6]) );
  NOR3_X1 U154 ( .A1(n619), .A2(n239), .A3(n629), .ZN(srl_result[7]) );
  NOR3_X1 U155 ( .A1(n420), .A2(n238), .A3(n8), .ZN(sll_result[25]) );
  OR2_X1 U156 ( .A1(n377), .A2(n217), .ZN(n470) );
  NAND2_X1 U157 ( .A1(n505), .A2(n210), .ZN(n529) );
  NAND2_X1 U158 ( .A1(n349), .A2(n210), .ZN(n366) );
  INV_X1 U159 ( .A(n429), .ZN(n270) );
  INV_X1 U160 ( .A(n582), .ZN(n304) );
  INV_X1 U161 ( .A(n573), .ZN(n301) );
  INV_X1 U162 ( .A(n393), .ZN(n277) );
  INV_X1 U163 ( .A(n399), .ZN(n275) );
  INV_X1 U164 ( .A(n422), .ZN(n273) );
  INV_X1 U165 ( .A(n342), .ZN(n290) );
  INV_X1 U166 ( .A(n354), .ZN(n289) );
  OR2_X1 U167 ( .A1(n338), .A2(n209), .ZN(n341) );
  INV_X1 U168 ( .A(n489), .ZN(n259) );
  INV_X1 U169 ( .A(n501), .ZN(n265) );
  INV_X1 U170 ( .A(n504), .ZN(n253) );
  INV_X1 U171 ( .A(n345), .ZN(n294) );
  INV_X1 U172 ( .A(n348), .ZN(n307) );
  INV_X1 U173 ( .A(n572), .ZN(n308) );
  INV_X1 U174 ( .A(n584), .ZN(n305) );
  NOR3_X1 U175 ( .A1(n319), .A2(n206), .A3(n51), .ZN(n148) );
  NOR3_X1 U176 ( .A1(n316), .A2(n211), .A3(n31), .ZN(n94) );
  NOR3_X1 U177 ( .A1(n313), .A2(n216), .A3(n51), .ZN(n79) );
  NOR3_X1 U178 ( .A1(n312), .A2(alu_src2[4]), .A3(n51), .ZN(n75) );
  NOR3_X1 U179 ( .A1(n309), .A2(n239), .A3(n51), .ZN(n71) );
  CLKBUF_X1 U181 ( .A(n52), .Z(n25) );
  CLKBUF_X1 U183 ( .A(n51), .Z(n31) );
  CLKBUF_X1 U184 ( .A(n51), .Z(n33) );
  CLKBUF_X1 U185 ( .A(n51), .Z(n32) );
  CLKBUF_X1 U190 ( .A(n51), .Z(n29) );
  INV_X1 U194 ( .A(alu_src2[3]), .ZN(n219) );
  INV_X1 U195 ( .A(n215), .ZN(n211) );
  OAI211_X1 U196 ( .C1(n1), .C2(n241), .A(n80), .B(n81), .ZN(alu_result[31])
         );
  AOI221_X1 U197 ( .B1(alu_src2[19]), .B2(n5), .C1(n42), .C2(n48), .A(n248), 
        .ZN(n81) );
  AOI22_X1 U198 ( .A1(srl_result[31]), .A2(n54), .B1(sll_result[31]), .B2(n16), 
        .ZN(n80) );
  INV_X1 U199 ( .A(n83), .ZN(n248) );
  NAND2_X1 U201 ( .A1(n197), .A2(n198), .ZN(alu_result[0]) );
  AOI222_X1 U202 ( .A1(adder_result[0]), .A2(n23), .B1(srl_result[0]), .B2(n54), .C1(sll_result[0]), .C2(n16), .ZN(n197) );
  AOI221_X1 U203 ( .B1(n44), .B2(n199), .C1(sra_result_0_), .C2(n48), .A(n200), 
        .ZN(n198) );
  AOI21_X1 U204 ( .B1(alu_src2[27]), .B2(n108), .A(n109), .ZN(n106) );
  AOI22_X1 U205 ( .A1(alu_src2[15]), .A2(n6), .B1(sra_result_27_), .B2(n48), 
        .ZN(n105) );
  AOI222_X1 U206 ( .A1(adder_result[27]), .A2(n22), .B1(srl_result[27]), .B2(
        n54), .C1(sll_result[27]), .C2(n17), .ZN(n107) );
  AOI21_X1 U207 ( .B1(alu_src2[28]), .B2(n103), .A(n104), .ZN(n101) );
  AOI22_X1 U208 ( .A1(alu_src2[16]), .A2(n6), .B1(sra_result_28_), .B2(n48), 
        .ZN(n100) );
  AOI222_X1 U209 ( .A1(adder_result[28]), .A2(n22), .B1(srl_result[28]), .B2(
        n54), .C1(sll_result[28]), .C2(n16), .ZN(n102) );
  AOI21_X1 U210 ( .B1(alu_src2[29]), .B2(n98), .A(n99), .ZN(n96) );
  AOI22_X1 U211 ( .A1(alu_src2[17]), .A2(n5), .B1(sra_result_29_), .B2(n48), 
        .ZN(n95) );
  AOI222_X1 U212 ( .A1(adder_result[29]), .A2(n22), .B1(srl_result[29]), .B2(
        n54), .C1(sll_result[29]), .C2(n16), .ZN(n97) );
  AOI21_X1 U213 ( .B1(alu_src2[30]), .B2(n89), .A(n90), .ZN(n87) );
  AOI22_X1 U268 ( .A1(alu_src2[18]), .A2(n4), .B1(sra_result_30_), .B2(n48), 
        .ZN(n86) );
  AOI222_X1 U269 ( .A1(adder_result[30]), .A2(n22), .B1(srl_result[30]), .B2(
        n54), .C1(sll_result[30]), .C2(n16), .ZN(n88) );
  AOI21_X1 U270 ( .B1(alu_src2[25]), .B2(n118), .A(n119), .ZN(n116) );
  AOI22_X1 U271 ( .A1(alu_src2[13]), .A2(n5), .B1(sra_result_25_), .B2(n48), 
        .ZN(n115) );
  AOI222_X1 U272 ( .A1(adder_result[25]), .A2(n23), .B1(srl_result[25]), .B2(
        n54), .C1(sll_result[25]), .C2(n17), .ZN(n117) );
  AOI21_X1 U273 ( .B1(alu_src2[26]), .B2(n113), .A(n114), .ZN(n111) );
  AOI22_X1 U274 ( .A1(alu_src2[14]), .A2(n4), .B1(sra_result_26_), .B2(n48), 
        .ZN(n110) );
  AOI222_X1 U275 ( .A1(adder_result[26]), .A2(n23), .B1(srl_result[26]), .B2(
        n54), .C1(sll_result[26]), .C2(n17), .ZN(n112) );
  AOI21_X1 U277 ( .B1(alu_src2[12]), .B2(n187), .A(n188), .ZN(n185) );
  AOI22_X1 U278 ( .A1(n44), .A2(n6), .B1(sra_result_12_), .B2(n48), .ZN(n184)
         );
  AOI222_X1 U279 ( .A1(adder_result[12]), .A2(n22), .B1(srl_result[12]), .B2(
        n54), .C1(sll_result[12]), .C2(n18), .ZN(n186) );
  AOI21_X1 U280 ( .B1(alu_src2[13]), .B2(n182), .A(n183), .ZN(n180) );
  AOI22_X1 U281 ( .A1(n206), .A2(n5), .B1(sra_result_13_), .B2(n48), .ZN(n179)
         );
  AOI222_X1 U282 ( .A1(adder_result[13]), .A2(n23), .B1(srl_result[13]), .B2(
        n54), .C1(sll_result[13]), .C2(n18), .ZN(n181) );
  AOI21_X1 U283 ( .B1(alu_src2[14]), .B2(n177), .A(n178), .ZN(n175) );
  AOI22_X1 U284 ( .A1(n211), .A2(n4), .B1(sra_result_14_), .B2(n48), .ZN(n174)
         );
  AOI222_X1 U285 ( .A1(adder_result[14]), .A2(n22), .B1(srl_result[14]), .B2(
        n54), .C1(sll_result[14]), .C2(n18), .ZN(n176) );
  AOI21_X1 U286 ( .B1(alu_src2[15]), .B2(n172), .A(n173), .ZN(n170) );
  AOI22_X1 U287 ( .A1(n6), .A2(n216), .B1(sra_result_15_), .B2(n48), .ZN(n169)
         );
  AOI222_X1 U288 ( .A1(adder_result[15]), .A2(n23), .B1(srl_result[15]), .B2(
        n54), .C1(sll_result[15]), .C2(n18), .ZN(n171) );
  AOI21_X1 U289 ( .B1(alu_src2[16]), .B2(n167), .A(n168), .ZN(n165) );
  AOI22_X1 U290 ( .A1(n4), .A2(alu_src2[4]), .B1(sra_result_16_), .B2(n48), 
        .ZN(n164) );
  AOI222_X1 U291 ( .A1(adder_result[16]), .A2(n23), .B1(srl_result[16]), .B2(
        n54), .C1(sll_result[16]), .C2(n18), .ZN(n166) );
  AOI21_X1 U292 ( .B1(alu_src2[17]), .B2(n162), .A(n163), .ZN(n160) );
  AOI22_X1 U293 ( .A1(n6), .A2(n237), .B1(sra_result_17_), .B2(n48), .ZN(n159)
         );
  AOI222_X1 U294 ( .A1(adder_result[17]), .A2(n23), .B1(srl_result[17]), .B2(
        n54), .C1(sll_result[17]), .C2(n18), .ZN(n161) );
  AOI21_X1 U295 ( .B1(alu_src2[18]), .B2(n157), .A(n158), .ZN(n155) );
  AOI22_X1 U296 ( .A1(n4), .A2(alu_src2[6]), .B1(sra_result_18_), .B2(n48), 
        .ZN(n154) );
  AOI222_X1 U297 ( .A1(adder_result[18]), .A2(n23), .B1(srl_result[18]), .B2(
        n54), .C1(sll_result[18]), .C2(n17), .ZN(n156) );
  AOI21_X1 U298 ( .B1(alu_src2[19]), .B2(n152), .A(n153), .ZN(n150) );
  AOI22_X1 U299 ( .A1(n5), .A2(alu_src2[7]), .B1(sra_result_19_), .B2(n48), 
        .ZN(n149) );
  AOI222_X1 U300 ( .A1(adder_result[19]), .A2(n23), .B1(srl_result[19]), .B2(
        n54), .C1(sll_result[19]), .C2(n17), .ZN(n151) );
  AOI21_X1 U301 ( .B1(alu_src2[20]), .B2(n143), .A(n144), .ZN(n141) );
  AOI22_X1 U302 ( .A1(n4), .A2(alu_src2[8]), .B1(sra_result_20_), .B2(n48), 
        .ZN(n140) );
  AOI222_X1 U303 ( .A1(adder_result[20]), .A2(n23), .B1(srl_result[20]), .B2(
        n54), .C1(sll_result[20]), .C2(n17), .ZN(n142) );
  AOI21_X1 U304 ( .B1(alu_src2[21]), .B2(n138), .A(n139), .ZN(n136) );
  AOI22_X1 U305 ( .A1(n5), .A2(alu_src2[9]), .B1(sra_result_21_), .B2(n48), 
        .ZN(n135) );
  AOI222_X1 U306 ( .A1(adder_result[21]), .A2(n23), .B1(srl_result[21]), .B2(
        n54), .C1(sll_result[21]), .C2(n17), .ZN(n137) );
  AOI21_X1 U307 ( .B1(alu_src2[22]), .B2(n133), .A(n134), .ZN(n131) );
  AOI22_X1 U308 ( .A1(alu_src2[10]), .A2(n4), .B1(sra_result_22_), .B2(n48), 
        .ZN(n130) );
  AOI222_X1 U309 ( .A1(adder_result[22]), .A2(n23), .B1(srl_result[22]), .B2(
        n54), .C1(sll_result[22]), .C2(n17), .ZN(n132) );
  AOI21_X1 U310 ( .B1(alu_src2[23]), .B2(n128), .A(n129), .ZN(n126) );
  AOI22_X1 U311 ( .A1(alu_src2[11]), .A2(n6), .B1(sra_result_23_), .B2(n48), 
        .ZN(n125) );
  AOI222_X1 U312 ( .A1(adder_result[23]), .A2(n23), .B1(srl_result[23]), .B2(
        n54), .C1(sll_result[23]), .C2(n17), .ZN(n127) );
  AOI21_X1 U313 ( .B1(alu_src2[24]), .B2(n123), .A(n124), .ZN(n121) );
  AOI22_X1 U314 ( .A1(alu_src2[12]), .A2(n5), .B1(sra_result_24_), .B2(n48), 
        .ZN(n120) );
  AOI222_X1 U315 ( .A1(adder_result[24]), .A2(n23), .B1(srl_result[24]), .B2(
        n54), .C1(sll_result[24]), .C2(n17), .ZN(n122) );
  NAND2_X1 U316 ( .A1(n189), .A2(n190), .ZN(alu_result[11]) );
  AOI221_X1 U317 ( .B1(sra_result_11_), .B2(n48), .C1(alu_src2[11]), .C2(n191), 
        .A(n192), .ZN(n190) );
  AOI222_X1 U318 ( .A1(adder_result[11]), .A2(n22), .B1(srl_result[11]), .B2(
        n54), .C1(sll_result[11]), .C2(n18), .ZN(n189) );
  OAI22_X1 U319 ( .A1(n52), .A2(n291), .B1(alu_src1[11]), .B2(n51), .ZN(n191)
         );
  INV_X1 U320 ( .A(alu_src1[8]), .ZN(n297) );
  INV_X1 U321 ( .A(alu_src1[9]), .ZN(n295) );
  NAND2_X1 U322 ( .A1(n193), .A2(n194), .ZN(alu_result[10]) );
  AOI221_X1 U323 ( .B1(sra_result_10_), .B2(n48), .C1(alu_src2[10]), .C2(n195), 
        .A(n196), .ZN(n194) );
  AOI222_X1 U324 ( .A1(adder_result[10]), .A2(n23), .B1(srl_result[10]), .B2(
        n54), .C1(sll_result[10]), .C2(n18), .ZN(n193) );
  OAI22_X1 U325 ( .A1(n52), .A2(n293), .B1(alu_src1[10]), .B2(n33), .ZN(n195)
         );
  NAND2_X1 U326 ( .A1(n76), .A2(n77), .ZN(alu_result[3]) );
  AOI222_X1 U327 ( .A1(adder_result[3]), .A2(n22), .B1(srl_result[3]), .B2(n54), .C1(sll_result[3]), .C2(n16), .ZN(n76) );
  AOI221_X1 U328 ( .B1(sra_result_3_), .B2(n48), .C1(n216), .C2(n78), .A(n79), 
        .ZN(n77) );
  NOR4_X1 U329 ( .A1(n235), .A2(n226), .A3(n476), .A4(n470), .ZN(sll_result[3]) );
  NAND2_X1 U330 ( .A1(n64), .A2(n65), .ZN(alu_result[6]) );
  AOI222_X1 U331 ( .A1(adder_result[6]), .A2(n22), .B1(srl_result[6]), .B2(n54), .C1(sll_result[6]), .C2(n16), .ZN(n64) );
  AOI221_X1 U332 ( .B1(sra_result_6_), .B2(n48), .C1(alu_src2[6]), .C2(n66), 
        .A(n67), .ZN(n65) );
  NOR4_X1 U333 ( .A1(n236), .A2(n225), .A3(n476), .A4(n473), .ZN(sll_result[6]) );
  NAND2_X1 U334 ( .A1(n60), .A2(n61), .ZN(alu_result[7]) );
  AOI221_X1 U335 ( .B1(sra_result_7_), .B2(n48), .C1(alu_src2[7]), .C2(n62), 
        .A(n63), .ZN(n61) );
  AOI222_X1 U336 ( .A1(adder_result[7]), .A2(n22), .B1(srl_result[7]), .B2(n54), .C1(sll_result[7]), .C2(n16), .ZN(n60) );
  NOR3_X1 U337 ( .A1(n302), .A2(alu_src2[7]), .A3(n29), .ZN(n63) );
  NAND2_X1 U338 ( .A1(n56), .A2(n57), .ZN(alu_result[8]) );
  AOI221_X1 U339 ( .B1(sra_result_8_), .B2(n48), .C1(alu_src2[8]), .C2(n58), 
        .A(n59), .ZN(n57) );
  AOI222_X1 U340 ( .A1(adder_result[8]), .A2(n22), .B1(srl_result[8]), .B2(n54), .C1(sll_result[8]), .C2(n16), .ZN(n56) );
  NOR3_X1 U341 ( .A1(n297), .A2(alu_src2[8]), .A3(n29), .ZN(n59) );
  NAND2_X1 U342 ( .A1(n46), .A2(n47), .ZN(alu_result[9]) );
  AOI221_X1 U343 ( .B1(sra_result_9_), .B2(n48), .C1(alu_src2[9]), .C2(n49), 
        .A(n50), .ZN(n47) );
  AOI222_X1 U344 ( .A1(adder_result[9]), .A2(n22), .B1(srl_result[9]), .B2(n54), .C1(sll_result[9]), .C2(n17), .ZN(n46) );
  NOR3_X1 U345 ( .A1(n295), .A2(alu_src2[9]), .A3(n29), .ZN(n50) );
  NOR4_X1 U346 ( .A1(n325), .A2(alu_src2[10]), .A3(alu_src2[12]), .A4(
        alu_src2[11]), .ZN(n332) );
  NOR4_X1 U347 ( .A1(n327), .A2(alu_src2[23]), .A3(alu_src2[25]), .A4(
        alu_src2[24]), .ZN(n330) );
  NOR4_X1 U348 ( .A1(n326), .A2(alu_src2[16]), .A3(alu_src2[18]), .A4(
        alu_src2[17]), .ZN(n331) );
  NOR4_X1 U349 ( .A1(n478), .A2(alu_src2[10]), .A3(alu_src2[12]), .A4(
        alu_src2[11]), .ZN(n485) );
  NOR4_X1 U350 ( .A1(n480), .A2(alu_src2[23]), .A3(alu_src2[25]), .A4(
        alu_src2[24]), .ZN(n483) );
  NOR4_X1 U351 ( .A1(n479), .A2(alu_src2[16]), .A3(alu_src2[18]), .A4(
        alu_src2[17]), .ZN(n484) );
  NOR4_X1 U352 ( .A1(n639), .A2(alu_src2[29]), .A3(alu_src2[31]), .A4(
        alu_src2[30]), .ZN(n640) );
  OR4_X1 U353 ( .A1(alu_src2[7]), .A2(alu_src2[6]), .A3(alu_src2[9]), .A4(
        alu_src2[8]), .ZN(n639) );
  NOR4_X1 U354 ( .A1(n328), .A2(alu_src2[29]), .A3(alu_src2[31]), .A4(
        alu_src2[30]), .ZN(n329) );
  OR4_X1 U355 ( .A1(alu_src2[7]), .A2(alu_src2[6]), .A3(alu_src2[9]), .A4(
        alu_src2[8]), .ZN(n328) );
  NOR4_X1 U356 ( .A1(n481), .A2(alu_src2[29]), .A3(alu_src2[31]), .A4(
        alu_src2[30]), .ZN(n482) );
  OR4_X1 U357 ( .A1(alu_src2[7]), .A2(alu_src2[6]), .A3(alu_src2[9]), .A4(
        alu_src2[8]), .ZN(n481) );
  INV_X1 U358 ( .A(n215), .ZN(n212) );
  INV_X1 U359 ( .A(n215), .ZN(n213) );
  INV_X1 U360 ( .A(n215), .ZN(n214) );
  AOI21_X1 U361 ( .B1(n84), .B2(alu_src2[31]), .A(n85), .ZN(n83) );
  NOR3_X1 U362 ( .A1(n51), .A2(alu_src2[31]), .A3(n43), .ZN(n85) );
  OAI22_X1 U363 ( .A1(n51), .A2(n40), .B1(n43), .B2(n52), .ZN(n84) );
  INV_X1 U364 ( .A(alu_src1[13]), .ZN(n285) );
  INV_X1 U365 ( .A(alu_src1[14]), .ZN(n284) );
  INV_X1 U366 ( .A(alu_src1[15]), .ZN(n283) );
  INV_X1 U367 ( .A(alu_src1[16]), .ZN(n282) );
  INV_X1 U368 ( .A(alu_src1[17]), .ZN(n281) );
  INV_X1 U369 ( .A(alu_src1[18]), .ZN(n280) );
  OR4_X1 U371 ( .A1(alu_src2[20]), .A2(alu_src2[19]), .A3(alu_src2[22]), .A4(
        alu_src2[21]), .ZN(n637) );
  OR4_X1 U372 ( .A1(alu_src2[20]), .A2(alu_src2[19]), .A3(alu_src2[22]), .A4(
        alu_src2[21]), .ZN(n326) );
  OR4_X1 U373 ( .A1(alu_src2[20]), .A2(alu_src2[19]), .A3(alu_src2[22]), .A4(
        alu_src2[21]), .ZN(n479) );
  NOR4_X1 U375 ( .A1(n636), .A2(alu_src2[10]), .A3(alu_src2[12]), .A4(
        alu_src2[11]), .ZN(n643) );
  NOR4_X1 U376 ( .A1(n638), .A2(alu_src2[23]), .A3(alu_src2[25]), .A4(
        alu_src2[24]), .ZN(n641) );
  NOR4_X1 U377 ( .A1(n637), .A2(alu_src2[16]), .A3(alu_src2[18]), .A4(
        alu_src2[17]), .ZN(n642) );
  INV_X1 U378 ( .A(alu_src1[19]), .ZN(n279) );
  INV_X1 U379 ( .A(alu_src1[12]), .ZN(n287) );
  INV_X1 U380 ( .A(alu_src1[21]), .ZN(n276) );
  INV_X1 U381 ( .A(alu_src1[20]), .ZN(n278) );
  INV_X1 U382 ( .A(alu_src1[10]), .ZN(n293) );
  INV_X1 U383 ( .A(alu_src1[11]), .ZN(n291) );
  INV_X1 U384 ( .A(alu_src1[7]), .ZN(n302) );
  INV_X1 U385 ( .A(alu_src1[22]), .ZN(n274) );
  OR3_X1 U386 ( .A1(alu_src2[28]), .A2(alu_src2[27]), .A3(alu_src2[26]), .ZN(
        n638) );
  OR3_X1 U387 ( .A1(alu_src2[15]), .A2(alu_src2[14]), .A3(alu_src2[13]), .ZN(
        n636) );
  OR3_X1 U388 ( .A1(alu_src2[28]), .A2(alu_src2[27]), .A3(alu_src2[26]), .ZN(
        n327) );
  OR3_X1 U389 ( .A1(alu_src2[15]), .A2(alu_src2[14]), .A3(alu_src2[13]), .ZN(
        n325) );
  OR3_X1 U390 ( .A1(alu_src2[28]), .A2(alu_src2[27]), .A3(alu_src2[26]), .ZN(
        n480) );
  OR3_X1 U391 ( .A1(alu_src2[15]), .A2(alu_src2[14]), .A3(alu_src2[13]), .ZN(
        n478) );
  NAND2_X1 U392 ( .A1(n355), .A2(n215), .ZN(n377) );
  NAND2_X1 U393 ( .A1(alu_src1[0]), .A2(n205), .ZN(n338) );
  INV_X1 U394 ( .A(n511), .ZN(n250) );
  INV_X1 U395 ( .A(n510), .ZN(n256) );
  INV_X1 U396 ( .A(n509), .ZN(n262) );
  INV_X1 U397 ( .A(n508), .ZN(n268) );
  INV_X1 U398 ( .A(n333), .ZN(n292) );
  INV_X1 U399 ( .A(n340), .ZN(n286) );
  INV_X1 U400 ( .A(n336), .ZN(n310) );
  INV_X1 U401 ( .A(n335), .ZN(n303) );
  INV_X1 U402 ( .A(n337), .ZN(n315) );
  INV_X1 U403 ( .A(n334), .ZN(n296) );
  INV_X1 U404 ( .A(n549), .ZN(n311) );
  NOR3_X1 U405 ( .A1(n306), .A2(alu_src2[6]), .A3(n29), .ZN(n67) );
  NOR3_X1 U406 ( .A1(n293), .A2(alu_src2[10]), .A3(n29), .ZN(n196) );
  NOR3_X1 U407 ( .A1(n291), .A2(alu_src2[11]), .A3(n29), .ZN(n192) );
  OAI22_X1 U408 ( .A1(n52), .A2(n287), .B1(alu_src1[12]), .B2(n33), .ZN(n187)
         );
  OAI22_X1 U409 ( .A1(n52), .A2(n285), .B1(alu_src1[13]), .B2(n33), .ZN(n182)
         );
  OAI22_X1 U410 ( .A1(n52), .A2(n284), .B1(alu_src1[14]), .B2(n33), .ZN(n177)
         );
  OAI22_X1 U411 ( .A1(n52), .A2(n283), .B1(alu_src1[15]), .B2(n33), .ZN(n172)
         );
  OAI22_X1 U412 ( .A1(n25), .A2(n282), .B1(alu_src1[16]), .B2(n33), .ZN(n167)
         );
  OAI22_X1 U413 ( .A1(n25), .A2(n281), .B1(alu_src1[17]), .B2(n33), .ZN(n162)
         );
  OAI22_X1 U414 ( .A1(n25), .A2(n280), .B1(alu_src1[18]), .B2(n33), .ZN(n157)
         );
  OAI22_X1 U415 ( .A1(n25), .A2(n279), .B1(alu_src1[19]), .B2(n33), .ZN(n152)
         );
  OAI22_X1 U416 ( .A1(n25), .A2(n278), .B1(alu_src1[20]), .B2(n33), .ZN(n143)
         );
  OAI22_X1 U417 ( .A1(n25), .A2(n276), .B1(alu_src1[21]), .B2(n32), .ZN(n138)
         );
  OAI22_X1 U418 ( .A1(n25), .A2(n274), .B1(alu_src1[22]), .B2(n33), .ZN(n133)
         );
  OAI22_X1 U419 ( .A1(n25), .A2(n272), .B1(alu_src1[23]), .B2(n32), .ZN(n128)
         );
  OAI22_X1 U420 ( .A1(n25), .A2(n269), .B1(alu_src1[24]), .B2(n32), .ZN(n123)
         );
  OAI22_X1 U421 ( .A1(n25), .A2(n266), .B1(alu_src1[25]), .B2(n32), .ZN(n118)
         );
  OAI22_X1 U422 ( .A1(n25), .A2(n263), .B1(alu_src1[26]), .B2(n32), .ZN(n113)
         );
  OAI22_X1 U423 ( .A1(n52), .A2(n260), .B1(alu_src1[27]), .B2(n32), .ZN(n108)
         );
  OAI22_X1 U424 ( .A1(n52), .A2(n257), .B1(alu_src1[28]), .B2(n32), .ZN(n103)
         );
  OAI22_X1 U425 ( .A1(n52), .A2(n254), .B1(alu_src1[29]), .B2(n32), .ZN(n98)
         );
  OAI22_X1 U426 ( .A1(n25), .A2(n251), .B1(alu_src1[30]), .B2(n32), .ZN(n89)
         );
  OAI22_X1 U427 ( .A1(n25), .A2(n319), .B1(alu_src1[1]), .B2(n33), .ZN(n147)
         );
  OAI22_X1 U428 ( .A1(n52), .A2(n316), .B1(alu_src1[2]), .B2(n32), .ZN(n93) );
  OAI22_X1 U429 ( .A1(n52), .A2(n313), .B1(alu_src1[3]), .B2(n31), .ZN(n78) );
  OAI22_X1 U430 ( .A1(n52), .A2(n312), .B1(alu_src1[4]), .B2(n31), .ZN(n74) );
  OAI22_X1 U431 ( .A1(n52), .A2(n309), .B1(alu_src1[5]), .B2(n32), .ZN(n70) );
  OAI22_X1 U432 ( .A1(n52), .A2(n306), .B1(alu_src1[6]), .B2(n31), .ZN(n66) );
  OAI22_X1 U433 ( .A1(n52), .A2(n302), .B1(alu_src1[7]), .B2(n31), .ZN(n62) );
  OAI22_X1 U434 ( .A1(n52), .A2(n297), .B1(alu_src1[8]), .B2(n31), .ZN(n58) );
  OAI22_X1 U435 ( .A1(n295), .A2(n52), .B1(alu_src1[9]), .B2(n31), .ZN(n49) );
  NOR3_X1 U436 ( .A1(n287), .A2(alu_src2[12]), .A3(n29), .ZN(n188) );
  NOR3_X1 U437 ( .A1(n282), .A2(alu_src2[16]), .A3(n51), .ZN(n168) );
  NOR3_X1 U438 ( .A1(n281), .A2(alu_src2[17]), .A3(n29), .ZN(n163) );
  NOR3_X1 U439 ( .A1(n280), .A2(alu_src2[18]), .A3(n51), .ZN(n158) );
  NOR3_X1 U440 ( .A1(n272), .A2(alu_src2[23]), .A3(n31), .ZN(n129) );
  NOR3_X1 U441 ( .A1(n269), .A2(alu_src2[24]), .A3(n51), .ZN(n124) );
  NOR3_X1 U442 ( .A1(n266), .A2(alu_src2[25]), .A3(n51), .ZN(n119) );
  NOR3_X1 U443 ( .A1(n254), .A2(alu_src2[29]), .A3(n51), .ZN(n99) );
  NOR3_X1 U444 ( .A1(n251), .A2(alu_src2[30]), .A3(n31), .ZN(n90) );
  NOR3_X1 U445 ( .A1(n285), .A2(alu_src2[13]), .A3(n29), .ZN(n183) );
  NOR3_X1 U446 ( .A1(n284), .A2(alu_src2[14]), .A3(n29), .ZN(n178) );
  NOR3_X1 U447 ( .A1(n283), .A2(alu_src2[15]), .A3(n29), .ZN(n173) );
  NOR3_X1 U448 ( .A1(n279), .A2(alu_src2[19]), .A3(n51), .ZN(n153) );
  NOR3_X1 U449 ( .A1(n278), .A2(alu_src2[20]), .A3(n29), .ZN(n144) );
  NOR3_X1 U450 ( .A1(n276), .A2(alu_src2[21]), .A3(n51), .ZN(n139) );
  NOR3_X1 U451 ( .A1(n274), .A2(alu_src2[22]), .A3(n51), .ZN(n134) );
  NOR3_X1 U452 ( .A1(n263), .A2(alu_src2[26]), .A3(n31), .ZN(n114) );
  NOR3_X1 U453 ( .A1(n260), .A2(alu_src2[27]), .A3(n31), .ZN(n109) );
  NOR3_X1 U454 ( .A1(n257), .A2(alu_src2[28]), .A3(n31), .ZN(n104) );
  OAI22_X1 U455 ( .A1(n52), .A2(n320), .B1(alu_src1[0]), .B2(n32), .ZN(n199)
         );
  INV_X1 U457 ( .A(alu_src1[3]), .ZN(n313) );
  INV_X1 U458 ( .A(alu_src1[4]), .ZN(n312) );
  INV_X1 U459 ( .A(alu_src1[5]), .ZN(n309) );
  INV_X1 U460 ( .A(alu_src1[6]), .ZN(n306) );
  INV_X1 U461 ( .A(alu_src1[23]), .ZN(n272) );
  INV_X1 U462 ( .A(alu_src1[24]), .ZN(n269) );
  INV_X1 U463 ( .A(alu_src1[25]), .ZN(n266) );
  INV_X1 U464 ( .A(alu_src1[26]), .ZN(n263) );
  INV_X1 U465 ( .A(alu_src1[27]), .ZN(n260) );
  INV_X1 U466 ( .A(alu_src1[28]), .ZN(n257) );
  INV_X1 U467 ( .A(alu_src1[29]), .ZN(n254) );
  INV_X1 U468 ( .A(alu_src1[30]), .ZN(n251) );
  INV_X1 U469 ( .A(alu_src1[1]), .ZN(n319) );
  INV_X1 U470 ( .A(alu_src1[2]), .ZN(n316) );
  INV_X1 U471 ( .A(alu_src1[0]), .ZN(n320) );
  CLKBUF_X1 U472 ( .A(n55), .Z(n16) );
  CLKBUF_X1 U473 ( .A(n55), .Z(n17) );
  INV_X1 U474 ( .A(n1), .ZN(n23) );
  INV_X1 U475 ( .A(n1), .ZN(n22) );
  CLKBUF_X1 U476 ( .A(n55), .Z(n18) );
  NAND2_X1 U484 ( .A1(n202), .A2(n323), .ZN(n201) );
  OAI22_X1 U485 ( .A1(alu_control[0]), .A2(n241), .B1(adder_cout), .B2(n324), 
        .ZN(n202) );
  INV_X1 U486 ( .A(alu_src2[2]), .ZN(n215) );
  NOR4_X1 U487 ( .A1(n321), .A2(alu_control[0]), .A3(alu_control[1]), .A4(
        alu_control[2]), .ZN(n55) );
  INV_X1 U488 ( .A(alu_control[3]), .ZN(n321) );
  INV_X1 U489 ( .A(alu_control[1]), .ZN(n323) );
  INV_X1 U490 ( .A(alu_control[2]), .ZN(n322) );
  NOR3_X1 U491 ( .A1(n323), .A2(alu_control[2]), .A3(n321), .ZN(n203) );
  OR3_X1 U492 ( .A1(alu_control[0]), .A2(alu_control[3]), .A3(n323), .ZN(n1)
         );
  INV_X1 U494 ( .A(alu_control[0]), .ZN(n324) );
  CLKBUF_X1 U495 ( .A(n2), .Z(n4) );
  NOR4_X1 U496 ( .A1(n322), .A2(n321), .A3(n323), .A4(alu_control[0]), .ZN(n2)
         );
  CLKBUF_X1 U497 ( .A(n3), .Z(n5) );
  NOR4_X1 U498 ( .A1(n322), .A2(n321), .A3(n323), .A4(alu_control[0]), .ZN(n3)
         );
  CLKBUF_X1 U499 ( .A(n82), .Z(n6) );
  NOR4_X1 U500 ( .A1(n322), .A2(n321), .A3(n323), .A4(alu_control[0]), .ZN(n82) );
  INV_X1 U501 ( .A(alu_src1[31]), .ZN(n43) );
  INV_X1 U502 ( .A(alu_src2[0]), .ZN(n205) );
  INV_X1 U503 ( .A(alu_src2[1]), .ZN(n210) );
  CLKBUF_X1 U505 ( .A(alu_src2[4]), .Z(n223) );
  CLKBUF_X1 U506 ( .A(alu_src2[4]), .Z(n224) );
  CLKBUF_X1 U507 ( .A(alu_src2[4]), .Z(n225) );
  CLKBUF_X1 U508 ( .A(alu_src2[4]), .Z(n226) );
  CLKBUF_X1 U509 ( .A(alu_src2[4]), .Z(n227) );
  MUX2_X1 U511 ( .A(alu_src1[10]), .B(alu_src1[9]), .S(n44), .Z(n333) );
  MUX2_X1 U512 ( .A(alu_src1[8]), .B(alu_src1[7]), .S(n53), .Z(n334) );
  MUX2_X1 U513 ( .A(n292), .B(n296), .S(n209), .Z(n350) );
  MUX2_X1 U514 ( .A(alu_src1[6]), .B(alu_src1[5]), .S(n204), .Z(n335) );
  MUX2_X1 U515 ( .A(alu_src1[4]), .B(alu_src1[3]), .S(alu_src2[0]), .Z(n336)
         );
  MUX2_X1 U516 ( .A(n303), .B(n310), .S(n208), .Z(n352) );
  MUX2_X1 U517 ( .A(n350), .B(n352), .S(n211), .Z(n371) );
  MUX2_X1 U518 ( .A(alu_src1[2]), .B(alu_src1[1]), .S(n204), .Z(n337) );
  MUX2_X1 U519 ( .A(n315), .B(n338), .S(n208), .Z(n351) );
  MUX2_X1 U520 ( .A(n371), .B(n314), .S(n218), .Z(n425) );
  MUX2_X1 U521 ( .A(alu_src1[11]), .B(alu_src1[10]), .S(n204), .Z(n342) );
  MUX2_X1 U522 ( .A(alu_src1[9]), .B(alu_src1[8]), .S(n53), .Z(n344) );
  MUX2_X1 U523 ( .A(n342), .B(n344), .S(n208), .Z(n354) );
  MUX2_X1 U524 ( .A(alu_src1[7]), .B(alu_src1[6]), .S(n204), .Z(n343) );
  MUX2_X1 U525 ( .A(alu_src1[5]), .B(alu_src1[4]), .S(n53), .Z(n347) );
  MUX2_X1 U526 ( .A(n343), .B(n347), .S(n209), .Z(n356) );
  MUX2_X1 U527 ( .A(n354), .B(n356), .S(n214), .Z(n339) );
  MUX2_X1 U528 ( .A(alu_src1[3]), .B(alu_src1[2]), .S(n53), .Z(n346) );
  MUX2_X1 U529 ( .A(alu_src1[1]), .B(alu_src1[0]), .S(n204), .Z(n349) );
  MUX2_X1 U530 ( .A(n346), .B(n349), .S(n208), .Z(n355) );
  MUX2_X1 U531 ( .A(n288), .B(n377), .S(n218), .Z(n432) );
  MUX2_X1 U532 ( .A(alu_src1[12]), .B(alu_src1[11]), .S(n45), .Z(n340) );
  MUX2_X1 U533 ( .A(n286), .B(n292), .S(n209), .Z(n358) );
  MUX2_X1 U534 ( .A(n296), .B(n303), .S(n209), .Z(n360) );
  MUX2_X1 U535 ( .A(n358), .B(n360), .S(n212), .Z(n383) );
  MUX2_X1 U536 ( .A(n310), .B(n315), .S(n209), .Z(n359) );
  MUX2_X1 U537 ( .A(n359), .B(n341), .S(n212), .Z(n384) );
  MUX2_X1 U538 ( .A(n383), .B(n384), .S(n216), .Z(n440) );
  MUX2_X1 U539 ( .A(n285), .B(n287), .S(n53), .Z(n353) );
  MUX2_X1 U540 ( .A(n353), .B(n290), .S(n209), .Z(n365) );
  MUX2_X1 U541 ( .A(n344), .B(n343), .S(n209), .Z(n345) );
  MUX2_X1 U542 ( .A(n365), .B(n294), .S(n213), .Z(n389) );
  MUX2_X1 U543 ( .A(n347), .B(n346), .S(n209), .Z(n348) );
  MUX2_X1 U544 ( .A(n307), .B(n366), .S(alu_src2[2]), .Z(n390) );
  MUX2_X1 U545 ( .A(n389), .B(n390), .S(n218), .Z(n448) );
  MUX2_X1 U546 ( .A(n284), .B(n285), .S(n204), .Z(n357) );
  MUX2_X1 U547 ( .A(n357), .B(n286), .S(n209), .Z(n370) );
  MUX2_X1 U548 ( .A(n370), .B(n350), .S(n214), .Z(n395) );
  MUX2_X1 U549 ( .A(n352), .B(n351), .S(n214), .Z(n396) );
  MUX2_X1 U550 ( .A(n395), .B(n396), .S(n218), .Z(n458) );
  MUX2_X1 U551 ( .A(n283), .B(n284), .S(n204), .Z(n364) );
  MUX2_X1 U552 ( .A(n364), .B(n353), .S(n209), .Z(n376) );
  MUX2_X1 U553 ( .A(n376), .B(n289), .S(n212), .Z(n401) );
  MUX2_X1 U554 ( .A(n356), .B(n355), .S(n213), .Z(n402) );
  MUX2_X1 U555 ( .A(n401), .B(n298), .S(alu_src2[3]), .Z(n467) );
  MUX2_X1 U556 ( .A(n282), .B(n283), .S(n204), .Z(n369) );
  MUX2_X1 U557 ( .A(n369), .B(n357), .S(n209), .Z(n382) );
  MUX2_X1 U558 ( .A(n382), .B(n358), .S(n212), .Z(n407) );
  MUX2_X1 U559 ( .A(n360), .B(n359), .S(n213), .Z(n410) );
  MUX2_X1 U560 ( .A(n407), .B(n410), .S(n217), .Z(n362) );
  MUX2_X1 U561 ( .A(n362), .B(n361), .S(n223), .Z(n363) );
  MUX2_X1 U562 ( .A(n281), .B(n282), .S(n204), .Z(n375) );
  MUX2_X1 U563 ( .A(n375), .B(n364), .S(n209), .Z(n388) );
  MUX2_X1 U564 ( .A(n388), .B(n365), .S(n213), .Z(n415) );
  MUX2_X1 U565 ( .A(n294), .B(n307), .S(n214), .Z(n418) );
  MUX2_X1 U566 ( .A(n415), .B(n418), .S(alu_src2[3]), .Z(n367) );
  MUX2_X1 U567 ( .A(n367), .B(n380), .S(n232), .Z(n368) );
  MUX2_X1 U568 ( .A(n280), .B(n281), .S(n204), .Z(n381) );
  MUX2_X1 U569 ( .A(n381), .B(n369), .S(n209), .Z(n394) );
  MUX2_X1 U570 ( .A(n394), .B(n370), .S(alu_src2[2]), .Z(n424) );
  MUX2_X1 U571 ( .A(n424), .B(n371), .S(alu_src2[3]), .Z(n373) );
  MUX2_X1 U572 ( .A(n373), .B(n451), .S(n232), .Z(n374) );
  MUX2_X1 U573 ( .A(n279), .B(n280), .S(n204), .Z(n387) );
  MUX2_X1 U574 ( .A(n387), .B(n375), .S(n209), .Z(n400) );
  MUX2_X1 U575 ( .A(n400), .B(n376), .S(alu_src2[2]), .Z(n431) );
  MUX2_X1 U576 ( .A(n431), .B(n288), .S(n217), .Z(n378) );
  MUX2_X1 U577 ( .A(n378), .B(n470), .S(n232), .Z(n379) );
  MUX2_X1 U578 ( .A(alu_src1[20]), .B(alu_src1[19]), .S(n204), .Z(n393) );
  MUX2_X1 U579 ( .A(n277), .B(n381), .S(n209), .Z(n406) );
  MUX2_X1 U580 ( .A(n406), .B(n382), .S(alu_src2[2]), .Z(n439) );
  MUX2_X1 U581 ( .A(n439), .B(n383), .S(n218), .Z(n385) );
  MUX2_X1 U582 ( .A(n385), .B(n471), .S(n232), .Z(n386) );
  MUX2_X1 U583 ( .A(alu_src1[21]), .B(alu_src1[20]), .S(n204), .Z(n399) );
  MUX2_X1 U584 ( .A(n275), .B(n387), .S(n209), .Z(n414) );
  MUX2_X1 U585 ( .A(n414), .B(n388), .S(alu_src2[2]), .Z(n447) );
  MUX2_X1 U586 ( .A(n447), .B(n389), .S(n218), .Z(n391) );
  MUX2_X1 U587 ( .A(n391), .B(n472), .S(n232), .Z(n392) );
  MUX2_X1 U588 ( .A(alu_src1[22]), .B(alu_src1[21]), .S(n204), .Z(n405) );
  MUX2_X1 U589 ( .A(n405), .B(n393), .S(n209), .Z(n422) );
  MUX2_X1 U590 ( .A(n273), .B(n394), .S(alu_src2[2]), .Z(n457) );
  MUX2_X1 U591 ( .A(n457), .B(n395), .S(n218), .Z(n397) );
  MUX2_X1 U592 ( .A(n397), .B(n473), .S(n232), .Z(n398) );
  MUX2_X1 U593 ( .A(alu_src1[23]), .B(alu_src1[22]), .S(n204), .Z(n413) );
  MUX2_X1 U594 ( .A(n413), .B(n399), .S(n209), .Z(n429) );
  MUX2_X1 U595 ( .A(n270), .B(n400), .S(n211), .Z(n466) );
  MUX2_X1 U596 ( .A(n466), .B(n401), .S(n218), .Z(n403) );
  MUX2_X1 U597 ( .A(n403), .B(n474), .S(n232), .Z(n404) );
  MUX2_X1 U598 ( .A(alu_src1[24]), .B(alu_src1[23]), .S(n204), .Z(n421) );
  MUX2_X1 U599 ( .A(n421), .B(n405), .S(n209), .Z(n436) );
  MUX2_X1 U600 ( .A(n267), .B(n406), .S(alu_src2[2]), .Z(n408) );
  MUX2_X1 U601 ( .A(n408), .B(n407), .S(n218), .Z(n411) );
  MUX2_X1 U602 ( .A(n410), .B(n317), .S(n218), .Z(n475) );
  MUX2_X1 U603 ( .A(n411), .B(n475), .S(n232), .Z(n412) );
  MUX2_X1 U604 ( .A(alu_src1[25]), .B(alu_src1[24]), .S(n204), .Z(n428) );
  MUX2_X1 U605 ( .A(n428), .B(n413), .S(n209), .Z(n444) );
  MUX2_X1 U606 ( .A(n264), .B(n414), .S(alu_src2[2]), .Z(n416) );
  MUX2_X1 U607 ( .A(n416), .B(n415), .S(n218), .Z(n419) );
  MUX2_X1 U608 ( .A(n418), .B(n318), .S(n218), .Z(n477) );
  MUX2_X1 U609 ( .A(n419), .B(n477), .S(n232), .Z(n420) );
  MUX2_X1 U610 ( .A(alu_src1[26]), .B(alu_src1[25]), .S(n204), .Z(n435) );
  MUX2_X1 U611 ( .A(n435), .B(n421), .S(n209), .Z(n454) );
  MUX2_X1 U612 ( .A(n454), .B(n422), .S(alu_src2[2]), .Z(n423) );
  MUX2_X1 U613 ( .A(n261), .B(n424), .S(n218), .Z(n426) );
  MUX2_X1 U614 ( .A(n426), .B(n425), .S(n232), .Z(n427) );
  MUX2_X1 U615 ( .A(alu_src1[27]), .B(alu_src1[26]), .S(n204), .Z(n443) );
  MUX2_X1 U616 ( .A(n443), .B(n428), .S(n208), .Z(n463) );
  MUX2_X1 U617 ( .A(n463), .B(n429), .S(alu_src2[2]), .Z(n430) );
  MUX2_X1 U618 ( .A(n258), .B(n431), .S(n218), .Z(n433) );
  MUX2_X1 U619 ( .A(n433), .B(n432), .S(n232), .Z(n434) );
  MUX2_X1 U620 ( .A(alu_src1[28]), .B(alu_src1[27]), .S(n204), .Z(n452) );
  MUX2_X1 U621 ( .A(n452), .B(n435), .S(n208), .Z(n437) );
  MUX2_X1 U622 ( .A(n437), .B(n436), .S(alu_src2[2]), .Z(n438) );
  MUX2_X1 U623 ( .A(n255), .B(n439), .S(n218), .Z(n441) );
  MUX2_X1 U624 ( .A(n441), .B(n440), .S(n232), .Z(n442) );
  MUX2_X1 U625 ( .A(alu_src1[29]), .B(alu_src1[28]), .S(n204), .Z(n461) );
  MUX2_X1 U626 ( .A(n461), .B(n443), .S(n208), .Z(n445) );
  MUX2_X1 U627 ( .A(n445), .B(n444), .S(alu_src2[2]), .Z(n446) );
  MUX2_X1 U628 ( .A(n252), .B(n447), .S(n218), .Z(n449) );
  MUX2_X1 U629 ( .A(n449), .B(n448), .S(n231), .Z(n450) );
  MUX2_X1 U630 ( .A(alu_src1[30]), .B(alu_src1[29]), .S(n204), .Z(n453) );
  MUX2_X1 U631 ( .A(n453), .B(n452), .S(n208), .Z(n455) );
  MUX2_X1 U632 ( .A(n455), .B(n454), .S(alu_src2[2]), .Z(n456) );
  MUX2_X1 U633 ( .A(n249), .B(n457), .S(n218), .Z(n459) );
  MUX2_X1 U634 ( .A(n459), .B(n458), .S(n231), .Z(n460) );
  MUX2_X1 U635 ( .A(n40), .B(alu_src1[30]), .S(n53), .Z(n462) );
  MUX2_X1 U636 ( .A(n462), .B(n461), .S(n208), .Z(n464) );
  MUX2_X1 U637 ( .A(n464), .B(n463), .S(alu_src2[2]), .Z(n465) );
  MUX2_X1 U638 ( .A(n466), .B(n242), .S(n219), .Z(n468) );
  MUX2_X1 U639 ( .A(n468), .B(n467), .S(n231), .Z(n469) );
  MUX2_X1 U641 ( .A(n297), .B(n295), .S(n53), .Z(n574) );
  MUX2_X1 U642 ( .A(n293), .B(n291), .S(n53), .Z(n494) );
  MUX2_X1 U643 ( .A(n574), .B(n494), .S(n208), .Z(n593) );
  MUX2_X1 U644 ( .A(n287), .B(n285), .S(n53), .Z(n493) );
  MUX2_X1 U645 ( .A(n284), .B(n283), .S(n53), .Z(n496) );
  MUX2_X1 U646 ( .A(n493), .B(n496), .S(n208), .Z(n515) );
  MUX2_X1 U647 ( .A(n593), .B(n515), .S(alu_src2[2]), .Z(n621) );
  MUX2_X1 U648 ( .A(alu_src1[0]), .B(alu_src1[1]), .S(n53), .Z(n486) );
  MUX2_X1 U649 ( .A(alu_src1[2]), .B(alu_src1[3]), .S(n53), .Z(n571) );
  MUX2_X1 U650 ( .A(n486), .B(n571), .S(n208), .Z(n487) );
  MUX2_X1 U651 ( .A(alu_src1[4]), .B(alu_src1[5]), .S(n53), .Z(n570) );
  MUX2_X1 U652 ( .A(alu_src1[6]), .B(alu_src1[7]), .S(n53), .Z(n573) );
  MUX2_X1 U653 ( .A(n570), .B(n573), .S(n208), .Z(n592) );
  MUX2_X1 U654 ( .A(n487), .B(n592), .S(alu_src2[2]), .Z(n488) );
  MUX2_X1 U655 ( .A(n621), .B(n299), .S(n219), .Z(n491) );
  MUX2_X1 U656 ( .A(n282), .B(n281), .S(n53), .Z(n495) );
  MUX2_X1 U657 ( .A(n280), .B(n279), .S(n53), .Z(n498) );
  MUX2_X1 U658 ( .A(n495), .B(n498), .S(n208), .Z(n514) );
  MUX2_X1 U659 ( .A(n278), .B(n276), .S(n53), .Z(n497) );
  MUX2_X1 U660 ( .A(alu_src1[22]), .B(alu_src1[23]), .S(n53), .Z(n500) );
  MUX2_X1 U661 ( .A(n497), .B(n271), .S(n208), .Z(n516) );
  MUX2_X1 U662 ( .A(n514), .B(n516), .S(alu_src2[2]), .Z(n620) );
  MUX2_X1 U663 ( .A(alu_src1[24]), .B(alu_src1[25]), .S(n53), .Z(n499) );
  MUX2_X1 U664 ( .A(alu_src1[26]), .B(alu_src1[27]), .S(n53), .Z(n503) );
  MUX2_X1 U665 ( .A(n499), .B(n503), .S(n208), .Z(n489) );
  MUX2_X1 U666 ( .A(alu_src1[28]), .B(alu_src1[29]), .S(n53), .Z(n502) );
  MUX2_X1 U667 ( .A(alu_src1[30]), .B(n40), .S(n53), .Z(n505) );
  MUX2_X1 U668 ( .A(n502), .B(n505), .S(n208), .Z(n490) );
  MUX2_X1 U669 ( .A(n259), .B(n244), .S(alu_src2[2]), .Z(n564) );
  MUX2_X1 U670 ( .A(n620), .B(n564), .S(n218), .Z(n539) );
  MUX2_X1 U671 ( .A(n491), .B(n539), .S(n231), .Z(n492) );
  MUX2_X1 U672 ( .A(n494), .B(n493), .S(n208), .Z(n606) );
  MUX2_X1 U673 ( .A(n496), .B(n495), .S(n208), .Z(n528) );
  MUX2_X1 U674 ( .A(n606), .B(n528), .S(n214), .Z(n575) );
  MUX2_X1 U675 ( .A(n498), .B(n497), .S(n208), .Z(n527) );
  MUX2_X1 U676 ( .A(n500), .B(n499), .S(n208), .Z(n501) );
  MUX2_X1 U677 ( .A(n527), .B(n265), .S(n214), .Z(n545) );
  MUX2_X1 U678 ( .A(n575), .B(n545), .S(n218), .Z(n506) );
  MUX2_X1 U679 ( .A(n503), .B(n502), .S(n208), .Z(n504) );
  MUX2_X1 U680 ( .A(n253), .B(n529), .S(n214), .Z(n544) );
  MUX2_X1 U681 ( .A(n506), .B(n566), .S(n231), .Z(n507) );
  MUX2_X1 U682 ( .A(n291), .B(n287), .S(n45), .Z(n550) );
  MUX2_X1 U683 ( .A(n285), .B(n284), .S(n45), .Z(n520) );
  MUX2_X1 U684 ( .A(n550), .B(n520), .S(n207), .Z(n613) );
  MUX2_X1 U685 ( .A(n283), .B(n282), .S(n45), .Z(n519) );
  MUX2_X1 U686 ( .A(n281), .B(n280), .S(n45), .Z(n522) );
  MUX2_X1 U687 ( .A(n519), .B(n522), .S(n207), .Z(n533) );
  MUX2_X1 U688 ( .A(n613), .B(n533), .S(n214), .Z(n587) );
  MUX2_X1 U689 ( .A(n279), .B(n278), .S(n45), .Z(n521) );
  MUX2_X1 U690 ( .A(n276), .B(n274), .S(n45), .Z(n523) );
  MUX2_X1 U691 ( .A(n521), .B(n523), .S(n207), .Z(n532) );
  MUX2_X1 U692 ( .A(alu_src1[23]), .B(alu_src1[24]), .S(n45), .Z(n508) );
  MUX2_X1 U693 ( .A(alu_src1[25]), .B(alu_src1[26]), .S(n45), .Z(n509) );
  MUX2_X1 U694 ( .A(n268), .B(n262), .S(n207), .Z(n535) );
  MUX2_X1 U695 ( .A(n532), .B(n535), .S(n214), .Z(n547) );
  MUX2_X1 U696 ( .A(n587), .B(n547), .S(n218), .Z(n512) );
  MUX2_X1 U697 ( .A(alu_src1[27]), .B(alu_src1[28]), .S(n45), .Z(n510) );
  MUX2_X1 U698 ( .A(alu_src1[29]), .B(alu_src1[30]), .S(n45), .Z(n511) );
  MUX2_X1 U699 ( .A(n256), .B(n250), .S(n207), .Z(n534) );
  MUX2_X1 U700 ( .A(n534), .B(n536), .S(n214), .Z(n546) );
  MUX2_X1 U701 ( .A(n512), .B(n567), .S(n231), .Z(n513) );
  MUX2_X1 U702 ( .A(n515), .B(n514), .S(n214), .Z(n594) );
  MUX2_X1 U703 ( .A(n516), .B(n259), .S(n214), .Z(n557) );
  MUX2_X1 U704 ( .A(n594), .B(n557), .S(n218), .Z(n517) );
  MUX2_X1 U705 ( .A(n517), .B(n568), .S(n231), .Z(n518) );
  MUX2_X1 U706 ( .A(n520), .B(n519), .S(n207), .Z(n551) );
  MUX2_X1 U707 ( .A(n522), .B(n521), .S(n207), .Z(n541) );
  MUX2_X1 U708 ( .A(n551), .B(n541), .S(n214), .Z(n601) );
  MUX2_X1 U709 ( .A(n523), .B(n268), .S(n207), .Z(n540) );
  MUX2_X1 U710 ( .A(n262), .B(n256), .S(n207), .Z(n543) );
  MUX2_X1 U711 ( .A(n540), .B(n543), .S(n214), .Z(n559) );
  MUX2_X1 U712 ( .A(n601), .B(n559), .S(n218), .Z(n525) );
  MUX2_X1 U713 ( .A(n250), .B(n524), .S(n207), .Z(n542) );
  MUX2_X1 U714 ( .A(n525), .B(n569), .S(n231), .Z(n526) );
  MUX2_X1 U715 ( .A(n528), .B(n527), .S(n214), .Z(n608) );
  MUX2_X1 U716 ( .A(n265), .B(n253), .S(n214), .Z(n561) );
  MUX2_X1 U717 ( .A(n608), .B(n561), .S(alu_src2[3]), .Z(n530) );
  MUX2_X1 U718 ( .A(n530), .B(n580), .S(n231), .Z(n531) );
  MUX2_X1 U719 ( .A(n533), .B(n532), .S(n214), .Z(n615) );
  MUX2_X1 U720 ( .A(n535), .B(n534), .S(n214), .Z(n563) );
  MUX2_X1 U721 ( .A(n615), .B(n563), .S(alu_src2[3]), .Z(n537) );
  MUX2_X1 U722 ( .A(n537), .B(n581), .S(n231), .Z(n538) );
  MUX2_X1 U723 ( .A(n541), .B(n540), .S(n214), .Z(n625) );
  MUX2_X1 U724 ( .A(n543), .B(n542), .S(n214), .Z(n565) );
  MUX2_X1 U725 ( .A(n625), .B(n565), .S(alu_src2[3]), .Z(n553) );
  MUX2_X1 U726 ( .A(n545), .B(n544), .S(alu_src2[3]), .Z(n577) );
  MUX2_X1 U727 ( .A(n547), .B(n546), .S(alu_src2[3]), .Z(n589) );
  MUX2_X1 U728 ( .A(alu_src1[1]), .B(alu_src1[2]), .S(n45), .Z(n548) );
  MUX2_X1 U729 ( .A(alu_src1[3]), .B(alu_src1[4]), .S(n45), .Z(n583) );
  MUX2_X1 U730 ( .A(n548), .B(n583), .S(n207), .Z(n549) );
  MUX2_X1 U731 ( .A(alu_src1[5]), .B(alu_src1[6]), .S(n45), .Z(n582) );
  MUX2_X1 U732 ( .A(n302), .B(n297), .S(n45), .Z(n586) );
  MUX2_X1 U733 ( .A(n304), .B(n586), .S(n207), .Z(n600) );
  MUX2_X1 U734 ( .A(n311), .B(n600), .S(n214), .Z(n552) );
  MUX2_X1 U735 ( .A(n295), .B(n293), .S(n45), .Z(n585) );
  MUX2_X1 U736 ( .A(n585), .B(n550), .S(n207), .Z(n599) );
  MUX2_X1 U737 ( .A(n599), .B(n551), .S(n213), .Z(n626) );
  MUX2_X1 U738 ( .A(n552), .B(n626), .S(alu_src2[3]), .Z(n554) );
  MUX2_X1 U739 ( .A(n554), .B(n553), .S(n231), .Z(n555) );
  MUX2_X1 U740 ( .A(n557), .B(n243), .S(alu_src2[3]), .Z(n596) );
  MUX2_X1 U741 ( .A(n559), .B(n247), .S(alu_src2[3]), .Z(n603) );
  MUX2_X1 U742 ( .A(n561), .B(n245), .S(alu_src2[3]), .Z(n610) );
  MUX2_X1 U743 ( .A(n563), .B(n246), .S(alu_src2[3]), .Z(n617) );
  MUX2_X1 U744 ( .A(n571), .B(n570), .S(n207), .Z(n572) );
  MUX2_X1 U745 ( .A(n301), .B(n574), .S(n207), .Z(n607) );
  MUX2_X1 U746 ( .A(n308), .B(n607), .S(n213), .Z(n576) );
  MUX2_X1 U747 ( .A(n576), .B(n575), .S(alu_src2[3]), .Z(n578) );
  MUX2_X1 U748 ( .A(n578), .B(n577), .S(n231), .Z(n579) );
  MUX2_X1 U749 ( .A(n583), .B(n582), .S(n207), .Z(n584) );
  MUX2_X1 U750 ( .A(n586), .B(n585), .S(n207), .Z(n614) );
  MUX2_X1 U751 ( .A(n305), .B(n614), .S(n213), .Z(n588) );
  MUX2_X1 U752 ( .A(n588), .B(n587), .S(alu_src2[3]), .Z(n590) );
  MUX2_X1 U753 ( .A(n590), .B(n589), .S(n231), .Z(n591) );
  MUX2_X1 U754 ( .A(n300), .B(n593), .S(n213), .Z(n595) );
  MUX2_X1 U755 ( .A(n595), .B(n594), .S(alu_src2[3]), .Z(n597) );
  MUX2_X1 U756 ( .A(n597), .B(n596), .S(n231), .Z(n598) );
  MUX2_X1 U757 ( .A(n600), .B(n599), .S(n213), .Z(n602) );
  MUX2_X1 U758 ( .A(n602), .B(n601), .S(alu_src2[3]), .Z(n604) );
  MUX2_X1 U759 ( .A(n604), .B(n603), .S(n230), .Z(n605) );
  MUX2_X1 U760 ( .A(n607), .B(n606), .S(n213), .Z(n609) );
  MUX2_X1 U761 ( .A(n609), .B(n608), .S(alu_src2[3]), .Z(n611) );
  MUX2_X1 U762 ( .A(n611), .B(n610), .S(n230), .Z(n612) );
  MUX2_X1 U763 ( .A(n614), .B(n613), .S(n213), .Z(n616) );
  MUX2_X1 U764 ( .A(n616), .B(n615), .S(alu_src2[3]), .Z(n618) );
  MUX2_X1 U765 ( .A(n618), .B(n617), .S(n230), .Z(n619) );
  MUX2_X1 U766 ( .A(n621), .B(n620), .S(alu_src2[3]), .Z(n623) );
  MUX2_X1 U767 ( .A(n623), .B(n622), .S(n230), .Z(n624) );
  MUX2_X1 U768 ( .A(n626), .B(n625), .S(n217), .Z(n628) );
  MUX2_X1 U769 ( .A(n628), .B(n627), .S(n230), .Z(n630) );
  MUX2_X1 U770 ( .A(alu_src1[0]), .B(alu_src1[1]), .S(n45), .Z(n631) );
  MUX2_X1 U771 ( .A(alu_src1[2]), .B(alu_src1[3]), .S(alu_src2[0]), .Z(n757)
         );
  MUX2_X1 U772 ( .A(n631), .B(n757), .S(alu_src2[1]), .Z(n632) );
  MUX2_X1 U773 ( .A(alu_src1[4]), .B(alu_src1[5]), .S(alu_src2[0]), .Z(n756)
         );
  MUX2_X1 U774 ( .A(alu_src1[6]), .B(alu_src1[7]), .S(alu_src2[0]), .Z(n759)
         );
  MUX2_X1 U775 ( .A(n756), .B(n759), .S(alu_src2[1]), .Z(n782) );
  MUX2_X1 U776 ( .A(n632), .B(n782), .S(n213), .Z(n633) );
  MUX2_X1 U777 ( .A(alu_src1[8]), .B(alu_src1[9]), .S(alu_src2[0]), .Z(n758)
         );
  MUX2_X1 U778 ( .A(alu_src1[10]), .B(alu_src1[11]), .S(alu_src2[0]), .Z(n646)
         );
  MUX2_X1 U779 ( .A(n758), .B(n646), .S(alu_src2[1]), .Z(n781) );
  MUX2_X1 U780 ( .A(alu_src1[12]), .B(alu_src1[13]), .S(alu_src2[0]), .Z(n645)
         );
  MUX2_X1 U781 ( .A(alu_src1[14]), .B(alu_src1[15]), .S(alu_src2[0]), .Z(n648)
         );
  MUX2_X1 U782 ( .A(n645), .B(n648), .S(alu_src2[1]), .Z(n663) );
  MUX2_X1 U783 ( .A(n781), .B(n663), .S(n213), .Z(n814) );
  MUX2_X1 U784 ( .A(n633), .B(n814), .S(n217), .Z(n634) );
  MUX2_X1 U785 ( .A(alu_src1[16]), .B(alu_src1[17]), .S(alu_src2[0]), .Z(n647)
         );
  MUX2_X1 U786 ( .A(alu_src1[18]), .B(alu_src1[19]), .S(alu_src2[0]), .Z(n650)
         );
  MUX2_X1 U787 ( .A(n647), .B(n650), .S(alu_src2[1]), .Z(n662) );
  MUX2_X1 U788 ( .A(alu_src1[20]), .B(alu_src1[21]), .S(n45), .Z(n649) );
  MUX2_X1 U789 ( .A(alu_src1[22]), .B(alu_src1[23]), .S(n44), .Z(n652) );
  MUX2_X1 U790 ( .A(n649), .B(n652), .S(alu_src2[1]), .Z(n665) );
  MUX2_X1 U791 ( .A(n662), .B(n665), .S(n213), .Z(n813) );
  MUX2_X1 U792 ( .A(alu_src1[24]), .B(alu_src1[25]), .S(n45), .Z(n651) );
  MUX2_X1 U793 ( .A(alu_src1[26]), .B(alu_src1[27]), .S(n45), .Z(n654) );
  MUX2_X1 U794 ( .A(n651), .B(n654), .S(n207), .Z(n664) );
  MUX2_X1 U795 ( .A(alu_src1[28]), .B(alu_src1[29]), .S(n45), .Z(n653) );
  MUX2_X1 U796 ( .A(alu_src1[30]), .B(alu_src1[31]), .S(n45), .Z(n655) );
  MUX2_X1 U797 ( .A(n653), .B(n655), .S(n206), .Z(n666) );
  MUX2_X1 U798 ( .A(n664), .B(n666), .S(n213), .Z(n738) );
  MUX2_X1 U799 ( .A(n813), .B(n738), .S(n217), .Z(n697) );
  MUX2_X1 U800 ( .A(n634), .B(n697), .S(n230), .Z(n635) );
  MUX2_X1 U801 ( .A(n635), .B(alu_src1[31]), .S(n239), .Z(n644) );
  MUX2_X1 U802 ( .A(n42), .B(n644), .S(n824), .Z(sra_result_0_) );
  MUX2_X1 U803 ( .A(n646), .B(n645), .S(alu_src2[1]), .Z(n797) );
  MUX2_X1 U804 ( .A(n648), .B(n647), .S(alu_src2[1]), .Z(n683) );
  MUX2_X1 U805 ( .A(n797), .B(n683), .S(n213), .Z(n761) );
  MUX2_X1 U806 ( .A(n650), .B(n649), .S(n207), .Z(n682) );
  MUX2_X1 U807 ( .A(n652), .B(n651), .S(n207), .Z(n685) );
  MUX2_X1 U808 ( .A(n682), .B(n685), .S(n213), .Z(n707) );
  MUX2_X1 U809 ( .A(n761), .B(n707), .S(n217), .Z(n656) );
  MUX2_X1 U810 ( .A(n654), .B(n653), .S(n207), .Z(n684) );
  MUX2_X1 U811 ( .A(n655), .B(n42), .S(n207), .Z(n686) );
  MUX2_X1 U812 ( .A(n684), .B(n686), .S(n213), .Z(n706) );
  MUX2_X1 U813 ( .A(n706), .B(alu_src1[31]), .S(n217), .Z(n744) );
  MUX2_X1 U814 ( .A(n656), .B(n744), .S(n230), .Z(n657) );
  MUX2_X1 U815 ( .A(n657), .B(alu_src1[31]), .S(n239), .Z(n658) );
  MUX2_X1 U816 ( .A(n41), .B(n658), .S(n824), .Z(sra_result_10_) );
  MUX2_X1 U817 ( .A(alu_src1[11]), .B(alu_src1[12]), .S(alu_src2[0]), .Z(n716)
         );
  MUX2_X1 U818 ( .A(alu_src1[13]), .B(alu_src1[14]), .S(alu_src2[0]), .Z(n671)
         );
  MUX2_X1 U819 ( .A(n716), .B(n671), .S(alu_src2[1]), .Z(n805) );
  MUX2_X1 U820 ( .A(alu_src1[15]), .B(alu_src1[16]), .S(alu_src2[0]), .Z(n670)
         );
  MUX2_X1 U821 ( .A(alu_src1[17]), .B(alu_src1[18]), .S(n44), .Z(n673) );
  MUX2_X1 U822 ( .A(n670), .B(n673), .S(alu_src2[1]), .Z(n691) );
  MUX2_X1 U823 ( .A(n805), .B(n691), .S(n213), .Z(n775) );
  MUX2_X1 U824 ( .A(alu_src1[19]), .B(alu_src1[20]), .S(n44), .Z(n672) );
  MUX2_X1 U825 ( .A(alu_src1[21]), .B(alu_src1[22]), .S(n44), .Z(n675) );
  MUX2_X1 U826 ( .A(n672), .B(n675), .S(alu_src2[1]), .Z(n690) );
  MUX2_X1 U827 ( .A(alu_src1[23]), .B(alu_src1[24]), .S(n44), .Z(n674) );
  MUX2_X1 U828 ( .A(alu_src1[25]), .B(alu_src1[26]), .S(n44), .Z(n677) );
  MUX2_X1 U829 ( .A(n674), .B(n677), .S(alu_src2[1]), .Z(n693) );
  MUX2_X1 U830 ( .A(n690), .B(n693), .S(n213), .Z(n711) );
  MUX2_X1 U831 ( .A(n775), .B(n711), .S(n217), .Z(n659) );
  MUX2_X1 U832 ( .A(alu_src1[27]), .B(alu_src1[28]), .S(n44), .Z(n676) );
  MUX2_X1 U833 ( .A(alu_src1[29]), .B(alu_src1[30]), .S(n44), .Z(n678) );
  MUX2_X1 U834 ( .A(n676), .B(n678), .S(alu_src2[1]), .Z(n692) );
  MUX2_X1 U835 ( .A(n692), .B(alu_src1[31]), .S(n213), .Z(n710) );
  MUX2_X1 U836 ( .A(n710), .B(alu_src1[31]), .S(n217), .Z(n747) );
  MUX2_X1 U837 ( .A(n659), .B(n747), .S(n230), .Z(n660) );
  MUX2_X1 U838 ( .A(n660), .B(n42), .S(n239), .Z(n661) );
  MUX2_X1 U839 ( .A(n40), .B(n661), .S(n824), .Z(sra_result_11_) );
  MUX2_X1 U840 ( .A(n663), .B(n662), .S(n214), .Z(n783) );
  MUX2_X1 U841 ( .A(n665), .B(n664), .S(n212), .Z(n724) );
  MUX2_X1 U842 ( .A(n783), .B(n724), .S(n217), .Z(n667) );
  MUX2_X1 U843 ( .A(n666), .B(n42), .S(n212), .Z(n723) );
  MUX2_X1 U844 ( .A(n723), .B(n42), .S(n217), .Z(n750) );
  MUX2_X1 U845 ( .A(n667), .B(n750), .S(n230), .Z(n668) );
  MUX2_X1 U846 ( .A(n668), .B(n42), .S(n239), .Z(n669) );
  MUX2_X1 U847 ( .A(n40), .B(n669), .S(n824), .Z(sra_result_12_) );
  MUX2_X1 U848 ( .A(n671), .B(n670), .S(n206), .Z(n717) );
  MUX2_X1 U849 ( .A(n673), .B(n672), .S(n206), .Z(n701) );
  MUX2_X1 U850 ( .A(n717), .B(n701), .S(n212), .Z(n791) );
  MUX2_X1 U851 ( .A(n675), .B(n674), .S(n206), .Z(n700) );
  MUX2_X1 U852 ( .A(n677), .B(n676), .S(n206), .Z(n703) );
  MUX2_X1 U853 ( .A(n700), .B(n703), .S(n212), .Z(n728) );
  MUX2_X1 U854 ( .A(n791), .B(n728), .S(n217), .Z(n679) );
  MUX2_X1 U855 ( .A(n678), .B(n42), .S(n206), .Z(n702) );
  MUX2_X1 U856 ( .A(n702), .B(n42), .S(n212), .Z(n727) );
  MUX2_X1 U857 ( .A(n727), .B(n42), .S(n217), .Z(n753) );
  MUX2_X1 U858 ( .A(n679), .B(n753), .S(n230), .Z(n680) );
  MUX2_X1 U859 ( .A(n680), .B(n42), .S(n239), .Z(n681) );
  MUX2_X1 U860 ( .A(n40), .B(n681), .S(n824), .Z(sra_result_13_) );
  MUX2_X1 U861 ( .A(n683), .B(n682), .S(n212), .Z(n799) );
  MUX2_X1 U862 ( .A(n685), .B(n684), .S(n212), .Z(n732) );
  MUX2_X1 U863 ( .A(n799), .B(n732), .S(n217), .Z(n687) );
  MUX2_X1 U864 ( .A(n686), .B(n42), .S(n212), .Z(n731) );
  MUX2_X1 U865 ( .A(n731), .B(n42), .S(n217), .Z(n767) );
  MUX2_X1 U866 ( .A(n687), .B(n767), .S(n230), .Z(n688) );
  MUX2_X1 U867 ( .A(n688), .B(n42), .S(n239), .Z(n689) );
  MUX2_X1 U868 ( .A(n40), .B(n689), .S(n824), .Z(sra_result_14_) );
  MUX2_X1 U869 ( .A(n691), .B(n690), .S(n212), .Z(n807) );
  MUX2_X1 U870 ( .A(n693), .B(n692), .S(n213), .Z(n735) );
  MUX2_X1 U871 ( .A(n807), .B(n735), .S(n216), .Z(n694) );
  MUX2_X1 U872 ( .A(n694), .B(n42), .S(n230), .Z(n695) );
  MUX2_X1 U873 ( .A(n695), .B(n42), .S(n239), .Z(n696) );
  MUX2_X1 U874 ( .A(n40), .B(n696), .S(n824), .Z(sra_result_15_) );
  MUX2_X1 U875 ( .A(n697), .B(n42), .S(n230), .Z(n698) );
  MUX2_X1 U876 ( .A(n698), .B(n42), .S(n239), .Z(n699) );
  MUX2_X1 U877 ( .A(n40), .B(n699), .S(n824), .Z(sra_result_16_) );
  MUX2_X1 U878 ( .A(n701), .B(n700), .S(n212), .Z(n819) );
  MUX2_X1 U879 ( .A(n703), .B(n702), .S(n212), .Z(n741) );
  MUX2_X1 U880 ( .A(n819), .B(n741), .S(n217), .Z(n719) );
  MUX2_X1 U881 ( .A(n719), .B(n42), .S(n229), .Z(n704) );
  MUX2_X1 U882 ( .A(n704), .B(n42), .S(n239), .Z(n705) );
  MUX2_X1 U883 ( .A(n40), .B(n705), .S(n824), .Z(sra_result_17_) );
  MUX2_X1 U884 ( .A(n707), .B(n706), .S(n217), .Z(n763) );
  MUX2_X1 U885 ( .A(n763), .B(n42), .S(n229), .Z(n708) );
  MUX2_X1 U886 ( .A(n708), .B(n42), .S(n239), .Z(n709) );
  MUX2_X1 U887 ( .A(n40), .B(n709), .S(n824), .Z(sra_result_18_) );
  MUX2_X1 U888 ( .A(n711), .B(n710), .S(n217), .Z(n777) );
  MUX2_X1 U889 ( .A(n777), .B(n42), .S(n230), .Z(n712) );
  MUX2_X1 U890 ( .A(n712), .B(n41), .S(n239), .Z(n713) );
  MUX2_X1 U891 ( .A(n40), .B(n713), .S(n824), .Z(sra_result_19_) );
  MUX2_X1 U892 ( .A(alu_src1[1]), .B(alu_src1[2]), .S(n44), .Z(n714) );
  MUX2_X1 U893 ( .A(alu_src1[3]), .B(alu_src1[4]), .S(n44), .Z(n771) );
  MUX2_X1 U894 ( .A(n714), .B(n771), .S(n206), .Z(n715) );
  MUX2_X1 U895 ( .A(alu_src1[5]), .B(alu_src1[6]), .S(n44), .Z(n770) );
  MUX2_X1 U896 ( .A(alu_src1[7]), .B(alu_src1[8]), .S(n44), .Z(n773) );
  MUX2_X1 U897 ( .A(n770), .B(n773), .S(n206), .Z(n790) );
  MUX2_X1 U898 ( .A(n715), .B(n790), .S(n212), .Z(n718) );
  MUX2_X1 U899 ( .A(alu_src1[9]), .B(alu_src1[10]), .S(n44), .Z(n772) );
  MUX2_X1 U900 ( .A(n772), .B(n716), .S(n206), .Z(n789) );
  MUX2_X1 U901 ( .A(n789), .B(n717), .S(n212), .Z(n820) );
  MUX2_X1 U902 ( .A(n718), .B(n820), .S(n217), .Z(n720) );
  MUX2_X1 U903 ( .A(n720), .B(n719), .S(n229), .Z(n721) );
  MUX2_X1 U904 ( .A(n721), .B(n41), .S(n239), .Z(n722) );
  MUX2_X1 U905 ( .A(n42), .B(n722), .S(n824), .Z(sra_result_1_) );
  MUX2_X1 U906 ( .A(n724), .B(n723), .S(n217), .Z(n785) );
  MUX2_X1 U907 ( .A(n785), .B(n41), .S(n229), .Z(n725) );
  MUX2_X1 U908 ( .A(n725), .B(n41), .S(n239), .Z(n726) );
  MUX2_X1 U909 ( .A(n40), .B(n726), .S(n824), .Z(sra_result_20_) );
  MUX2_X1 U910 ( .A(n728), .B(n727), .S(n216), .Z(n793) );
  MUX2_X1 U911 ( .A(n793), .B(n41), .S(n229), .Z(n729) );
  MUX2_X1 U912 ( .A(n729), .B(n41), .S(n239), .Z(n730) );
  MUX2_X1 U913 ( .A(n42), .B(n730), .S(n824), .Z(sra_result_21_) );
  MUX2_X1 U914 ( .A(n732), .B(n731), .S(n216), .Z(n801) );
  MUX2_X1 U915 ( .A(n801), .B(n41), .S(n229), .Z(n733) );
  MUX2_X1 U916 ( .A(n733), .B(n41), .S(n239), .Z(n734) );
  MUX2_X1 U917 ( .A(n40), .B(n734), .S(n824), .Z(sra_result_22_) );
  MUX2_X1 U918 ( .A(n735), .B(n41), .S(n216), .Z(n809) );
  MUX2_X1 U919 ( .A(n809), .B(n41), .S(n229), .Z(n736) );
  MUX2_X1 U920 ( .A(n736), .B(n41), .S(n239), .Z(n737) );
  MUX2_X1 U921 ( .A(n40), .B(n737), .S(n824), .Z(sra_result_23_) );
  MUX2_X1 U922 ( .A(n738), .B(n41), .S(n216), .Z(n815) );
  MUX2_X1 U923 ( .A(n815), .B(n41), .S(n229), .Z(n739) );
  MUX2_X1 U924 ( .A(n739), .B(n41), .S(n239), .Z(n740) );
  MUX2_X1 U925 ( .A(n42), .B(n740), .S(n824), .Z(sra_result_24_) );
  MUX2_X1 U926 ( .A(n741), .B(n41), .S(n216), .Z(n821) );
  MUX2_X1 U927 ( .A(n821), .B(n41), .S(n229), .Z(n742) );
  MUX2_X1 U928 ( .A(n742), .B(n41), .S(n239), .Z(n743) );
  MUX2_X1 U929 ( .A(n42), .B(n743), .S(n824), .Z(sra_result_25_) );
  MUX2_X1 U930 ( .A(n744), .B(n41), .S(n229), .Z(n745) );
  MUX2_X1 U931 ( .A(n745), .B(n40), .S(n239), .Z(n746) );
  MUX2_X1 U932 ( .A(n40), .B(n746), .S(n824), .Z(sra_result_26_) );
  MUX2_X1 U933 ( .A(n747), .B(n41), .S(n229), .Z(n748) );
  MUX2_X1 U934 ( .A(n748), .B(n42), .S(alu_src2[5]), .Z(n749) );
  MUX2_X1 U935 ( .A(n40), .B(n749), .S(n824), .Z(sra_result_27_) );
  MUX2_X1 U936 ( .A(n750), .B(n41), .S(n229), .Z(n751) );
  MUX2_X1 U937 ( .A(n751), .B(n41), .S(alu_src2[5]), .Z(n752) );
  MUX2_X1 U938 ( .A(n40), .B(n752), .S(n824), .Z(sra_result_28_) );
  MUX2_X1 U939 ( .A(n753), .B(n41), .S(n229), .Z(n754) );
  MUX2_X1 U940 ( .A(n754), .B(n41), .S(alu_src2[5]), .Z(n755) );
  MUX2_X1 U941 ( .A(n40), .B(n755), .S(n824), .Z(sra_result_29_) );
  MUX2_X1 U942 ( .A(n757), .B(n756), .S(n206), .Z(n760) );
  MUX2_X1 U943 ( .A(n759), .B(n758), .S(n206), .Z(n798) );
  MUX2_X1 U944 ( .A(n760), .B(n798), .S(n212), .Z(n762) );
  MUX2_X1 U945 ( .A(n762), .B(n761), .S(n216), .Z(n764) );
  MUX2_X1 U946 ( .A(n764), .B(n763), .S(n229), .Z(n765) );
  MUX2_X1 U947 ( .A(n765), .B(n41), .S(alu_src2[5]), .Z(n766) );
  MUX2_X1 U948 ( .A(n40), .B(n766), .S(n824), .Z(sra_result_2_) );
  MUX2_X1 U949 ( .A(n767), .B(n41), .S(alu_src2[4]), .Z(n768) );
  MUX2_X1 U950 ( .A(n768), .B(n40), .S(alu_src2[5]), .Z(n769) );
  MUX2_X1 U951 ( .A(n40), .B(n769), .S(n824), .Z(sra_result_30_) );
  MUX2_X1 U952 ( .A(n771), .B(n770), .S(n206), .Z(n774) );
  MUX2_X1 U953 ( .A(n773), .B(n772), .S(n206), .Z(n806) );
  MUX2_X1 U954 ( .A(n774), .B(n806), .S(n212), .Z(n776) );
  MUX2_X1 U955 ( .A(n776), .B(n775), .S(n216), .Z(n778) );
  MUX2_X1 U956 ( .A(n778), .B(n777), .S(alu_src2[4]), .Z(n779) );
  MUX2_X1 U957 ( .A(n779), .B(n41), .S(alu_src2[5]), .Z(n780) );
  MUX2_X1 U958 ( .A(n40), .B(n780), .S(n824), .Z(sra_result_3_) );
  MUX2_X1 U959 ( .A(n782), .B(n781), .S(n212), .Z(n784) );
  MUX2_X1 U960 ( .A(n784), .B(n783), .S(n216), .Z(n786) );
  MUX2_X1 U961 ( .A(n786), .B(n785), .S(alu_src2[4]), .Z(n787) );
  MUX2_X1 U962 ( .A(n787), .B(n40), .S(alu_src2[5]), .Z(n788) );
  MUX2_X1 U963 ( .A(n40), .B(n788), .S(n824), .Z(sra_result_4_) );
  MUX2_X1 U964 ( .A(n790), .B(n789), .S(n212), .Z(n792) );
  MUX2_X1 U965 ( .A(n792), .B(n791), .S(n216), .Z(n794) );
  MUX2_X1 U966 ( .A(n794), .B(n793), .S(alu_src2[4]), .Z(n795) );
  MUX2_X1 U967 ( .A(n795), .B(n40), .S(alu_src2[5]), .Z(n796) );
  MUX2_X1 U968 ( .A(n40), .B(n796), .S(n824), .Z(sra_result_5_) );
  MUX2_X1 U969 ( .A(n798), .B(n797), .S(n211), .Z(n800) );
  MUX2_X1 U970 ( .A(n800), .B(n799), .S(n216), .Z(n802) );
  MUX2_X1 U971 ( .A(n802), .B(n801), .S(n226), .Z(n803) );
  MUX2_X1 U972 ( .A(n803), .B(n40), .S(alu_src2[5]), .Z(n804) );
  MUX2_X1 U973 ( .A(n40), .B(n804), .S(n824), .Z(sra_result_6_) );
  MUX2_X1 U974 ( .A(n806), .B(n805), .S(n212), .Z(n808) );
  MUX2_X1 U975 ( .A(n808), .B(n807), .S(n216), .Z(n810) );
  MUX2_X1 U976 ( .A(n810), .B(n809), .S(n227), .Z(n811) );
  MUX2_X1 U977 ( .A(n811), .B(n41), .S(alu_src2[5]), .Z(n812) );
  MUX2_X1 U978 ( .A(n42), .B(n812), .S(n824), .Z(sra_result_7_) );
  MUX2_X1 U979 ( .A(n814), .B(n813), .S(n216), .Z(n816) );
  MUX2_X1 U980 ( .A(n816), .B(n815), .S(n224), .Z(n817) );
  MUX2_X1 U981 ( .A(n817), .B(n40), .S(alu_src2[5]), .Z(n818) );
  MUX2_X1 U982 ( .A(n40), .B(n818), .S(n824), .Z(sra_result_8_) );
  MUX2_X1 U983 ( .A(n820), .B(n819), .S(n216), .Z(n822) );
  MUX2_X1 U984 ( .A(n822), .B(n821), .S(n225), .Z(n823) );
  MUX2_X1 U985 ( .A(n823), .B(n40), .S(alu_src2[5]), .Z(n825) );
  MUX2_X1 U986 ( .A(n41), .B(n825), .S(n824), .Z(sra_result_9_) );
  AND2_X2 U4 ( .A1(n324), .A2(n203), .ZN(n54) );
  AND2_X2 U5 ( .A1(alu_control[0]), .A2(n203), .ZN(n48) );
  AND4_X2 U134 ( .A1(n642), .A2(n640), .A3(n641), .A4(n643), .ZN(n824) );
  NAND3_X1 U136 ( .A1(n322), .A2(n321), .A3(n323), .ZN(n52) );
  NAND4_X1 U137 ( .A1(n485), .A2(n483), .A3(n482), .A4(n484), .ZN(n629) );
  NAND4_X1 U138 ( .A1(n332), .A2(n330), .A3(n329), .A4(n331), .ZN(n476) );
  NAND3_X1 U139 ( .A1(n322), .A2(n321), .A3(alu_control[0]), .ZN(n51) );
  NAND2_X2 U148 ( .A1(n22), .A2(n322), .ZN(N96) );
endmodule


module alu_control ( instr_30, func3, ALUOP, ALU_control );
  input [2:0] func3;
  input [1:0] ALUOP;
  output [3:0] ALU_control;
  input instr_30;
  wire   N42, N43, N44, N45, N46, n7, n8, n9, n10, n11, n12, n1, n2, n3, n4,
         n5, n6;

  DLH_X1 ALU_control_reg_3_ ( .G(N42), .D(N46), .Q(ALU_control[3]) );
  DLH_X1 ALU_control_reg_2_ ( .G(N42), .D(N45), .Q(ALU_control[2]) );
  DLH_X1 ALU_control_reg_1_ ( .G(N42), .D(N44), .Q(ALU_control[1]) );
  DLH_X1 ALU_control_reg_0_ ( .G(N42), .D(N43), .Q(ALU_control[0]) );
  NAND4_X1 U19 ( .A1(instr_30), .A2(n6), .A3(n4), .A4(n2), .ZN(n8) );
  AOI21_X1 U3 ( .B1(n2), .B2(func3[1]), .A(n5), .ZN(n7) );
  OAI211_X1 U4 ( .C1(func3[1]), .C2(n4), .A(n6), .B(n5), .ZN(N42) );
  OAI22_X1 U5 ( .A1(ALUOP[1]), .A2(ALUOP[0]), .B1(n10), .B2(n5), .ZN(N43) );
  AOI22_X1 U6 ( .A1(n11), .A2(func3[0]), .B1(func3[2]), .B2(n1), .ZN(n10) );
  INV_X1 U7 ( .A(n12), .ZN(n1) );
  NOR2_X1 U8 ( .A1(func3[2]), .A2(n3), .ZN(n11) );
  AOI21_X1 U9 ( .B1(n3), .B2(instr_30), .A(n4), .ZN(n12) );
  INV_X1 U10 ( .A(func3[0]), .ZN(n4) );
  INV_X1 U11 ( .A(ALUOP[1]), .ZN(n5) );
  INV_X1 U12 ( .A(func3[1]), .ZN(n3) );
  OAI21_X1 U13 ( .B1(func3[1]), .B2(n4), .A(n7), .ZN(N46) );
  INV_X1 U14 ( .A(ALUOP[0]), .ZN(n6) );
  INV_X1 U15 ( .A(func3[2]), .ZN(n2) );
  NAND2_X1 U16 ( .A1(n7), .A2(n8), .ZN(N45) );
  NAND2_X1 U17 ( .A1(ALUOP[1]), .A2(n9), .ZN(N44) );
  OAI21_X1 U18 ( .B1(func3[2]), .B2(n4), .A(n3), .ZN(n9) );
endmodule


module REG_WB ( clk, wdata, wa, regwrite, memtoreg, wdata_WB, wa_WB, 
        regwrite_WB, memtoreg_WB );
  input [31:0] wdata;
  input [4:0] wa;
  output [31:0] wdata_WB;
  output [4:0] wa_WB;
  input clk, regwrite, memtoreg;
  output regwrite_WB, memtoreg_WB;


  DFF_X1 wdata_WB_reg_31_ ( .D(wdata[31]), .CK(clk), .Q(wdata_WB[31]) );
  DFF_X1 wdata_WB_reg_30_ ( .D(wdata[30]), .CK(clk), .Q(wdata_WB[30]) );
  DFF_X1 wdata_WB_reg_29_ ( .D(wdata[29]), .CK(clk), .Q(wdata_WB[29]) );
  DFF_X1 wdata_WB_reg_28_ ( .D(wdata[28]), .CK(clk), .Q(wdata_WB[28]) );
  DFF_X1 wdata_WB_reg_27_ ( .D(wdata[27]), .CK(clk), .Q(wdata_WB[27]) );
  DFF_X1 wdata_WB_reg_26_ ( .D(wdata[26]), .CK(clk), .Q(wdata_WB[26]) );
  DFF_X1 wdata_WB_reg_25_ ( .D(wdata[25]), .CK(clk), .Q(wdata_WB[25]) );
  DFF_X1 wdata_WB_reg_24_ ( .D(wdata[24]), .CK(clk), .Q(wdata_WB[24]) );
  DFF_X1 wdata_WB_reg_23_ ( .D(wdata[23]), .CK(clk), .Q(wdata_WB[23]) );
  DFF_X1 wdata_WB_reg_22_ ( .D(wdata[22]), .CK(clk), .Q(wdata_WB[22]) );
  DFF_X1 wdata_WB_reg_21_ ( .D(wdata[21]), .CK(clk), .Q(wdata_WB[21]) );
  DFF_X1 wdata_WB_reg_20_ ( .D(wdata[20]), .CK(clk), .Q(wdata_WB[20]) );
  DFF_X1 wdata_WB_reg_19_ ( .D(wdata[19]), .CK(clk), .Q(wdata_WB[19]) );
  DFF_X1 wdata_WB_reg_18_ ( .D(wdata[18]), .CK(clk), .Q(wdata_WB[18]) );
  DFF_X1 wdata_WB_reg_17_ ( .D(wdata[17]), .CK(clk), .Q(wdata_WB[17]) );
  DFF_X1 wdata_WB_reg_16_ ( .D(wdata[16]), .CK(clk), .Q(wdata_WB[16]) );
  DFF_X1 wdata_WB_reg_15_ ( .D(wdata[15]), .CK(clk), .Q(wdata_WB[15]) );
  DFF_X1 wdata_WB_reg_14_ ( .D(wdata[14]), .CK(clk), .Q(wdata_WB[14]) );
  DFF_X1 wdata_WB_reg_13_ ( .D(wdata[13]), .CK(clk), .Q(wdata_WB[13]) );
  DFF_X1 wdata_WB_reg_12_ ( .D(wdata[12]), .CK(clk), .Q(wdata_WB[12]) );
  DFF_X1 wdata_WB_reg_11_ ( .D(wdata[11]), .CK(clk), .Q(wdata_WB[11]) );
  DFF_X1 wdata_WB_reg_10_ ( .D(wdata[10]), .CK(clk), .Q(wdata_WB[10]) );
  DFF_X1 wdata_WB_reg_9_ ( .D(wdata[9]), .CK(clk), .Q(wdata_WB[9]) );
  DFF_X1 wdata_WB_reg_8_ ( .D(wdata[8]), .CK(clk), .Q(wdata_WB[8]) );
  DFF_X1 wdata_WB_reg_7_ ( .D(wdata[7]), .CK(clk), .Q(wdata_WB[7]) );
  DFF_X1 wdata_WB_reg_6_ ( .D(wdata[6]), .CK(clk), .Q(wdata_WB[6]) );
  DFF_X1 wdata_WB_reg_5_ ( .D(wdata[5]), .CK(clk), .Q(wdata_WB[5]) );
  DFF_X1 wdata_WB_reg_4_ ( .D(wdata[4]), .CK(clk), .Q(wdata_WB[4]) );
  DFF_X1 wdata_WB_reg_3_ ( .D(wdata[3]), .CK(clk), .Q(wdata_WB[3]) );
  DFF_X1 wdata_WB_reg_2_ ( .D(wdata[2]), .CK(clk), .Q(wdata_WB[2]) );
  DFF_X1 wdata_WB_reg_1_ ( .D(wdata[1]), .CK(clk), .Q(wdata_WB[1]) );
  DFF_X1 wdata_WB_reg_0_ ( .D(wdata[0]), .CK(clk), .Q(wdata_WB[0]) );
  DFF_X1 wa_WB_reg_4_ ( .D(wa[4]), .CK(clk), .Q(wa_WB[4]) );
  DFF_X1 wa_WB_reg_3_ ( .D(wa[3]), .CK(clk), .Q(wa_WB[3]) );
  DFF_X1 wa_WB_reg_2_ ( .D(wa[2]), .CK(clk), .Q(wa_WB[2]) );
  DFF_X1 wa_WB_reg_1_ ( .D(wa[1]), .CK(clk), .Q(wa_WB[1]) );
  DFF_X1 wa_WB_reg_0_ ( .D(wa[0]), .CK(clk), .Q(wa_WB[0]) );
  DFF_X1 regwrite_WB_reg ( .D(regwrite), .CK(clk), .Q(regwrite_WB) );
endmodule


module Forward ( regwrite_WB, wa_WB, ra1_EX, ra2_EX, forwardA, forwardB );
  input [4:0] wa_WB;
  input [4:0] ra1_EX;
  input [4:0] ra2_EX;
  input regwrite_WB;
  output forwardA, forwardB;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  XOR2_X1 U9 ( .A(wa_WB[4]), .B(ra2_EX[4]), .Z(n4) );
  XOR2_X1 U10 ( .A(wa_WB[1]), .B(ra2_EX[1]), .Z(n3) );
  XOR2_X1 U11 ( .A(wa_WB[3]), .B(ra2_EX[3]), .Z(n2) );
  NAND4_X1 U12 ( .A1(n5), .A2(n6), .A3(regwrite_WB), .A4(n7), .ZN(n1) );
  XOR2_X1 U13 ( .A(wa_WB[1]), .B(ra1_EX[1]), .Z(n11) );
  XOR2_X1 U14 ( .A(wa_WB[4]), .B(ra1_EX[4]), .Z(n10) );
  XOR2_X1 U15 ( .A(wa_WB[3]), .B(ra1_EX[3]), .Z(n9) );
  NAND4_X1 U16 ( .A1(n12), .A2(n13), .A3(regwrite_WB), .A4(n7), .ZN(n8) );
  NOR4_X1 U1 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(forwardB) );
  XNOR2_X1 U2 ( .A(wa_WB[0]), .B(ra2_EX[0]), .ZN(n6) );
  XNOR2_X1 U3 ( .A(wa_WB[2]), .B(ra2_EX[2]), .ZN(n5) );
  XNOR2_X1 U4 ( .A(wa_WB[0]), .B(ra1_EX[0]), .ZN(n13) );
  XNOR2_X1 U5 ( .A(wa_WB[2]), .B(ra1_EX[2]), .ZN(n12) );
  OR4_X1 U6 ( .A1(wa_WB[3]), .A2(wa_WB[4]), .A3(wa_WB[2]), .A4(n14), .ZN(n7)
         );
  OR2_X1 U7 ( .A1(wa_WB[1]), .A2(wa_WB[0]), .ZN(n14) );
  NOR4_X1 U8 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(forwardA) );
endmodule


module RISC_V ( in, clk, alu_output_data );
  input [31:0] in;
  output [31:0] alu_output_data;
  input clk;
  wire   instr_6, instr_5, instr_4, instr_3, instr_2, instr_1, instr_0,
         regwrite_WB, ALUsrc, regwrite, funct7_EX, ALUsrc_EX, regwrite_EX,
         forwardA, forwardB, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n137, n139, n140, n148, n151, n153;
  wire   [4:0] wa;
  wire   [31:25] instr;
  wire   [2:0] funct3;
  wire   [4:0] ra1;
  wire   [4:0] ra2;
  wire   [4:0] wa_WB;
  wire   [31:0] rda;
  wire   [31:0] rdb;
  wire   [31:0] imm;
  wire   [1:0] ALUOP;
  wire   [31:0] rda_EX;
  wire   [31:0] rdb_EX;
  wire   [31:0] imm_EX;
  wire   [2:0] funct3_EX;
  wire   [4:0] wa_EX;
  wire   [1:0] ALUOP_EX;
  wire   [4:0] ra1_EX;
  wire   [4:0] ra2_EX;
  wire   [3:0] operation;
  wire   [31:0] alu_result;

  REG_ID REG_ID ( .clk(clk), .in(in), .instr({instr, ra2, ra1, funct3, wa, 
        instr_6, instr_5, instr_4, instr_3, instr_2, instr_1, instr_0}) );
  regfile regfile ( .clk(clk), .ra1(ra1), .ra2(ra2), .en_write(regwrite_WB), 
        .wa(wa_WB), .wdata(alu_output_data), .rd1(rda), .rd2(rdb) );
  ImmGen ImmGen ( .instr({instr, ra2, ra1, funct3, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, instr_6, instr_5, instr_4, instr_3, instr_2, instr_1, instr_0}), 
        .imm_out(imm) );
  control control ( .opcode({instr_6, instr_5, instr_4, instr_3, instr_2, 
        instr_1, instr_0}), .ALUsrc(ALUsrc), .ALUOP(ALUOP), .regwrite(regwrite) );
  REG_EX REG_EX ( .clk(clk), .rda(rda), .rdb(rdb), .imm(imm), .wa(wa), 
        .funct7(instr[30]), .funct3(funct3), .ALUsrc(ALUsrc), .ALUOP(ALUOP), 
        .regwrite(regwrite), .branch(1'b0), .memread(1'b0), .memwrite(1'b0), 
        .memtoreg(1'b0), .ra1(ra1), .ra2(ra2), .rda_EX(rda_EX), .rdb_EX(rdb_EX), .imm_EX(imm_EX), .wa_EX(wa_EX), .funct7_EX(funct7_EX), .funct3_EX(funct3_EX), 
        .ALUsrc_EX(ALUsrc_EX), .ALUOP_EX(ALUOP_EX), .regwrite_EX(regwrite_EX), 
        .ra1_EX(ra1_EX), .ra2_EX(ra2_EX) );
  alu_32bit alu_32bit ( .alu_src1({n64, n63, n62, n61, n60, n59, n58, n57, n56, 
        n55, n54, n53, n52, n51, n50, n49, n48, n47, n46, n45, n44, n43, n42, 
        n41, n40, n39, n38, n37, n36, n35, n34, n33}), .alu_src2({n8, n9, n11, 
        n12, n13, n14, n15, n16, n17, n18, n19, n20, n22, n23, n24, n25, n26, 
        n27, n28, n29, n30, n31, n1, n2, n3, n4, n5, n6, n7, n10, n21, n32}), 
        .alu_control(operation), .alu_result(alu_result) );
  alu_control alu_control ( .instr_30(funct7_EX), .func3(funct3_EX), .ALUOP(
        ALUOP_EX), .ALU_control(operation) );
  REG_WB REG_WB ( .clk(clk), .wdata(alu_result), .wa(wa_EX), .regwrite(
        regwrite_EX), .memtoreg(1'b0), .wdata_WB(alu_output_data), .wa_WB(
        wa_WB), .regwrite_WB(regwrite_WB) );
  Forward Forward ( .regwrite_WB(regwrite_WB), .wa_WB(wa_WB), .ra1_EX(ra1_EX), 
        .ra2_EX(ra2_EX), .forwardA(forwardA), .forwardB(forwardB) );
  CLKBUF_X1 U134 ( .A(n68), .Z(n137) );
  INV_X1 U135 ( .A(n148), .ZN(n139) );
  INV_X1 U140 ( .A(n148), .ZN(n140) );
  INV_X1 U151 ( .A(n71), .ZN(n3) );
  AOI222_X1 U152 ( .A1(imm_EX[7]), .A2(ALUsrc_EX), .B1(rdb_EX[7]), .B2(n68), 
        .C1(alu_output_data[7]), .C2(n69), .ZN(n71) );
  INV_X1 U153 ( .A(n107), .ZN(n36) );
  AOI22_X1 U154 ( .A1(n148), .A2(rda_EX[3]), .B1(alu_output_data[3]), .B2(n139), .ZN(n107) );
  INV_X1 U155 ( .A(n78), .ZN(n10) );
  AOI222_X1 U156 ( .A1(imm_EX[2]), .A2(ALUsrc_EX), .B1(rdb_EX[2]), .B2(n137), 
        .C1(alu_output_data[2]), .C2(n69), .ZN(n78) );
  INV_X1 U157 ( .A(n132), .ZN(n33) );
  AOI22_X1 U158 ( .A1(n148), .A2(rda_EX[0]), .B1(alu_output_data[0]), .B2(n139), .ZN(n132) );
  INV_X1 U159 ( .A(n75), .ZN(n7) );
  AOI222_X1 U160 ( .A1(imm_EX[3]), .A2(ALUsrc_EX), .B1(rdb_EX[3]), .B2(n68), 
        .C1(alu_output_data[3]), .C2(n69), .ZN(n75) );
  INV_X1 U161 ( .A(n100), .ZN(n32) );
  AOI222_X1 U162 ( .A1(imm_EX[0]), .A2(ALUsrc_EX), .B1(rdb_EX[0]), .B2(n68), 
        .C1(alu_output_data[0]), .C2(n69), .ZN(n100) );
  INV_X1 U163 ( .A(n89), .ZN(n21) );
  AOI222_X1 U164 ( .A1(imm_EX[1]), .A2(ALUsrc_EX), .B1(rdb_EX[1]), .B2(n68), 
        .C1(alu_output_data[1]), .C2(n69), .ZN(n89) );
  INV_X1 U166 ( .A(n74), .ZN(n6) );
  AOI222_X1 U167 ( .A1(imm_EX[4]), .A2(ALUsrc_EX), .B1(rdb_EX[4]), .B2(n68), 
        .C1(alu_output_data[4]), .C2(n69), .ZN(n74) );
  INV_X1 U168 ( .A(n73), .ZN(n5) );
  AOI222_X1 U169 ( .A1(imm_EX[5]), .A2(ALUsrc_EX), .B1(rdb_EX[5]), .B2(n68), 
        .C1(alu_output_data[5]), .C2(n69), .ZN(n73) );
  INV_X1 U170 ( .A(n98), .ZN(n30) );
  AOI222_X1 U171 ( .A1(imm_EX[11]), .A2(n151), .B1(rdb_EX[11]), .B2(n68), .C1(
        alu_output_data[11]), .C2(n69), .ZN(n98) );
  INV_X1 U172 ( .A(n93), .ZN(n25) );
  AOI222_X1 U173 ( .A1(imm_EX[16]), .A2(n151), .B1(rdb_EX[16]), .B2(n68), .C1(
        alu_output_data[16]), .C2(n69), .ZN(n93) );
  INV_X1 U174 ( .A(n99), .ZN(n31) );
  AOI222_X1 U175 ( .A1(imm_EX[10]), .A2(n151), .B1(rdb_EX[10]), .B2(n68), .C1(
        alu_output_data[10]), .C2(n69), .ZN(n99) );
  INV_X1 U176 ( .A(n97), .ZN(n29) );
  AOI222_X1 U177 ( .A1(imm_EX[12]), .A2(n151), .B1(rdb_EX[12]), .B2(n68), .C1(
        alu_output_data[12]), .C2(n69), .ZN(n97) );
  INV_X1 U178 ( .A(n91), .ZN(n23) );
  AOI222_X1 U179 ( .A1(imm_EX[18]), .A2(n151), .B1(rdb_EX[18]), .B2(n68), .C1(
        alu_output_data[18]), .C2(n69), .ZN(n91) );
  INV_X1 U180 ( .A(n83), .ZN(n15) );
  AOI222_X1 U181 ( .A1(imm_EX[25]), .A2(ALUsrc_EX), .B1(rdb_EX[25]), .B2(n137), 
        .C1(alu_output_data[25]), .C2(n69), .ZN(n83) );
  INV_X1 U182 ( .A(n121), .ZN(n34) );
  AOI22_X1 U183 ( .A1(n148), .A2(rda_EX[1]), .B1(alu_output_data[1]), .B2(n139), .ZN(n121) );
  INV_X1 U184 ( .A(n129), .ZN(n45) );
  AOI22_X1 U185 ( .A1(n148), .A2(rda_EX[12]), .B1(alu_output_data[12]), .B2(
        n139), .ZN(n129) );
  INV_X1 U186 ( .A(n128), .ZN(n46) );
  AOI22_X1 U187 ( .A1(n148), .A2(rda_EX[13]), .B1(alu_output_data[13]), .B2(
        n139), .ZN(n128) );
  INV_X1 U188 ( .A(n127), .ZN(n47) );
  AOI22_X1 U189 ( .A1(n148), .A2(rda_EX[14]), .B1(alu_output_data[14]), .B2(
        n139), .ZN(n127) );
  INV_X1 U190 ( .A(n110), .ZN(n35) );
  AOI22_X1 U191 ( .A1(n148), .A2(rda_EX[2]), .B1(alu_output_data[2]), .B2(n140), .ZN(n110) );
  INV_X1 U192 ( .A(n70), .ZN(n2) );
  AOI222_X1 U193 ( .A1(imm_EX[8]), .A2(ALUsrc_EX), .B1(rdb_EX[8]), .B2(n68), 
        .C1(alu_output_data[8]), .C2(n69), .ZN(n70) );
  INV_X1 U194 ( .A(n67), .ZN(n1) );
  AOI222_X1 U195 ( .A1(imm_EX[9]), .A2(ALUsrc_EX), .B1(rdb_EX[9]), .B2(n68), 
        .C1(alu_output_data[9]), .C2(n69), .ZN(n67) );
  INV_X1 U196 ( .A(n72), .ZN(n4) );
  AOI222_X1 U197 ( .A1(imm_EX[6]), .A2(ALUsrc_EX), .B1(rdb_EX[6]), .B2(n68), 
        .C1(alu_output_data[6]), .C2(n69), .ZN(n72) );
  INV_X1 U198 ( .A(n96), .ZN(n28) );
  AOI222_X1 U199 ( .A1(imm_EX[13]), .A2(n151), .B1(rdb_EX[13]), .B2(n68), .C1(
        alu_output_data[13]), .C2(n69), .ZN(n96) );
  INV_X1 U200 ( .A(n90), .ZN(n22) );
  AOI222_X1 U201 ( .A1(imm_EX[19]), .A2(n151), .B1(rdb_EX[19]), .B2(n68), .C1(
        alu_output_data[19]), .C2(n69), .ZN(n90) );
  INV_X1 U202 ( .A(n95), .ZN(n27) );
  AOI222_X1 U203 ( .A1(imm_EX[14]), .A2(n151), .B1(rdb_EX[14]), .B2(n68), .C1(
        alu_output_data[14]), .C2(n69), .ZN(n95) );
  INV_X1 U204 ( .A(n104), .ZN(n39) );
  AOI22_X1 U205 ( .A1(n148), .A2(rda_EX[6]), .B1(alu_output_data[6]), .B2(n140), .ZN(n104) );
  INV_X1 U206 ( .A(n106), .ZN(n37) );
  AOI22_X1 U207 ( .A1(n148), .A2(rda_EX[4]), .B1(alu_output_data[4]), .B2(n140), .ZN(n106) );
  INV_X1 U208 ( .A(n105), .ZN(n38) );
  AOI22_X1 U209 ( .A1(n148), .A2(rda_EX[5]), .B1(alu_output_data[5]), .B2(n140), .ZN(n105) );
  INV_X1 U210 ( .A(n94), .ZN(n26) );
  AOI222_X1 U211 ( .A1(imm_EX[15]), .A2(n151), .B1(rdb_EX[15]), .B2(n68), .C1(
        alu_output_data[15]), .C2(n69), .ZN(n94) );
  INV_X1 U212 ( .A(n103), .ZN(n40) );
  AOI22_X1 U213 ( .A1(n148), .A2(rda_EX[7]), .B1(alu_output_data[7]), .B2(n140), .ZN(n103) );
  INV_X1 U214 ( .A(n102), .ZN(n41) );
  AOI22_X1 U215 ( .A1(n148), .A2(rda_EX[8]), .B1(alu_output_data[8]), .B2(n140), .ZN(n102) );
  INV_X1 U216 ( .A(n101), .ZN(n42) );
  AOI22_X1 U217 ( .A1(n148), .A2(rda_EX[9]), .B1(alu_output_data[9]), .B2(n140), .ZN(n101) );
  INV_X1 U218 ( .A(n131), .ZN(n43) );
  AOI22_X1 U219 ( .A1(n148), .A2(rda_EX[10]), .B1(alu_output_data[10]), .B2(
        n139), .ZN(n131) );
  INV_X1 U220 ( .A(n130), .ZN(n44) );
  AOI22_X1 U221 ( .A1(n148), .A2(rda_EX[11]), .B1(alu_output_data[11]), .B2(
        n139), .ZN(n130) );
  INV_X1 U222 ( .A(n88), .ZN(n20) );
  AOI222_X1 U223 ( .A1(imm_EX[20]), .A2(ALUsrc_EX), .B1(rdb_EX[20]), .B2(n137), 
        .C1(alu_output_data[20]), .C2(n69), .ZN(n88) );
  INV_X1 U224 ( .A(n122), .ZN(n52) );
  AOI22_X1 U225 ( .A1(n148), .A2(rda_EX[19]), .B1(alu_output_data[19]), .B2(
        n139), .ZN(n122) );
  INV_X1 U227 ( .A(n123), .ZN(n51) );
  AOI22_X1 U228 ( .A1(n148), .A2(rda_EX[18]), .B1(alu_output_data[18]), .B2(
        n139), .ZN(n123) );
  INV_X1 U230 ( .A(n92), .ZN(n24) );
  AOI222_X1 U231 ( .A1(imm_EX[17]), .A2(n151), .B1(rdb_EX[17]), .B2(n68), .C1(
        alu_output_data[17]), .C2(n69), .ZN(n92) );
  INV_X1 U232 ( .A(n85), .ZN(n17) );
  AOI222_X1 U233 ( .A1(imm_EX[23]), .A2(ALUsrc_EX), .B1(rdb_EX[23]), .B2(n137), 
        .C1(alu_output_data[23]), .C2(n69), .ZN(n85) );
  INV_X1 U234 ( .A(n79), .ZN(n11) );
  AOI222_X1 U235 ( .A1(imm_EX[29]), .A2(ALUsrc_EX), .B1(rdb_EX[29]), .B2(n137), 
        .C1(alu_output_data[29]), .C2(n69), .ZN(n79) );
  INV_X1 U236 ( .A(n84), .ZN(n16) );
  AOI222_X1 U237 ( .A1(imm_EX[24]), .A2(ALUsrc_EX), .B1(rdb_EX[24]), .B2(n137), 
        .C1(alu_output_data[24]), .C2(n69), .ZN(n84) );
  INV_X1 U238 ( .A(n77), .ZN(n9) );
  AOI222_X1 U239 ( .A1(imm_EX[30]), .A2(ALUsrc_EX), .B1(rdb_EX[30]), .B2(n137), 
        .C1(alu_output_data[30]), .C2(n69), .ZN(n77) );
  INV_X1 U240 ( .A(n124), .ZN(n50) );
  AOI22_X1 U241 ( .A1(n148), .A2(rda_EX[17]), .B1(alu_output_data[17]), .B2(
        n139), .ZN(n124) );
  INV_X1 U242 ( .A(n126), .ZN(n48) );
  AOI22_X1 U243 ( .A1(n148), .A2(rda_EX[15]), .B1(alu_output_data[15]), .B2(
        n139), .ZN(n126) );
  INV_X1 U244 ( .A(n118), .ZN(n55) );
  AOI22_X1 U245 ( .A1(n148), .A2(rda_EX[22]), .B1(alu_output_data[22]), .B2(
        n140), .ZN(n118) );
  INV_X1 U246 ( .A(n117), .ZN(n56) );
  AOI22_X1 U247 ( .A1(n148), .A2(rda_EX[23]), .B1(alu_output_data[23]), .B2(
        n140), .ZN(n117) );
  INV_X1 U248 ( .A(n115), .ZN(n58) );
  AOI22_X1 U249 ( .A1(n148), .A2(rda_EX[25]), .B1(alu_output_data[25]), .B2(
        n140), .ZN(n115) );
  INV_X1 U250 ( .A(n114), .ZN(n59) );
  AOI22_X1 U251 ( .A1(n148), .A2(rda_EX[26]), .B1(alu_output_data[26]), .B2(
        n140), .ZN(n114) );
  INV_X1 U252 ( .A(n113), .ZN(n60) );
  AOI22_X1 U253 ( .A1(n148), .A2(rda_EX[27]), .B1(alu_output_data[27]), .B2(
        n140), .ZN(n113) );
  INV_X1 U254 ( .A(n112), .ZN(n61) );
  AOI22_X1 U255 ( .A1(n148), .A2(rda_EX[28]), .B1(alu_output_data[28]), .B2(
        n140), .ZN(n112) );
  INV_X1 U256 ( .A(n109), .ZN(n63) );
  AOI22_X1 U257 ( .A1(n148), .A2(rda_EX[30]), .B1(alu_output_data[30]), .B2(
        n140), .ZN(n109) );
  INV_X1 U258 ( .A(n116), .ZN(n57) );
  AOI22_X1 U259 ( .A1(n148), .A2(rda_EX[24]), .B1(alu_output_data[24]), .B2(
        n140), .ZN(n116) );
  INV_X1 U260 ( .A(n111), .ZN(n62) );
  AOI22_X1 U261 ( .A1(n148), .A2(rda_EX[29]), .B1(alu_output_data[29]), .B2(
        n140), .ZN(n111) );
  INV_X1 U262 ( .A(n87), .ZN(n19) );
  AOI222_X1 U263 ( .A1(imm_EX[21]), .A2(ALUsrc_EX), .B1(rdb_EX[21]), .B2(n137), 
        .C1(alu_output_data[21]), .C2(n69), .ZN(n87) );
  INV_X1 U264 ( .A(n120), .ZN(n53) );
  AOI22_X1 U265 ( .A1(n148), .A2(rda_EX[20]), .B1(alu_output_data[20]), .B2(
        n140), .ZN(n120) );
  INV_X1 U266 ( .A(n119), .ZN(n54) );
  AOI22_X1 U267 ( .A1(n148), .A2(rda_EX[21]), .B1(alu_output_data[21]), .B2(
        n140), .ZN(n119) );
  INV_X1 U268 ( .A(n86), .ZN(n18) );
  AOI222_X1 U269 ( .A1(imm_EX[22]), .A2(ALUsrc_EX), .B1(rdb_EX[22]), .B2(n137), 
        .C1(alu_output_data[22]), .C2(n69), .ZN(n86) );
  INV_X1 U270 ( .A(n82), .ZN(n14) );
  AOI222_X1 U271 ( .A1(imm_EX[26]), .A2(ALUsrc_EX), .B1(rdb_EX[26]), .B2(n137), 
        .C1(alu_output_data[26]), .C2(n69), .ZN(n82) );
  INV_X1 U272 ( .A(n81), .ZN(n13) );
  AOI222_X1 U273 ( .A1(imm_EX[27]), .A2(ALUsrc_EX), .B1(rdb_EX[27]), .B2(n137), 
        .C1(alu_output_data[27]), .C2(n69), .ZN(n81) );
  INV_X1 U274 ( .A(n80), .ZN(n12) );
  AOI222_X1 U275 ( .A1(imm_EX[28]), .A2(ALUsrc_EX), .B1(rdb_EX[28]), .B2(n137), 
        .C1(alu_output_data[28]), .C2(n69), .ZN(n80) );
  INV_X1 U276 ( .A(n125), .ZN(n49) );
  AOI22_X1 U277 ( .A1(n148), .A2(rda_EX[16]), .B1(alu_output_data[16]), .B2(
        n139), .ZN(n125) );
  CLKBUF_X1 U278 ( .A(ALUsrc_EX), .Z(n151) );
  INV_X1 U279 ( .A(n108), .ZN(n64) );
  AOI22_X1 U280 ( .A1(n148), .A2(rda_EX[31]), .B1(alu_output_data[31]), .B2(
        n140), .ZN(n108) );
  INV_X1 U281 ( .A(n76), .ZN(n8) );
  AOI222_X1 U282 ( .A1(imm_EX[31]), .A2(ALUsrc_EX), .B1(rdb_EX[31]), .B2(n68), 
        .C1(alu_output_data[31]), .C2(n69), .ZN(n76) );
  INV_X2 U133 ( .A(forwardA), .ZN(n148) );
  AND2_X2 U136 ( .A1(n153), .A2(forwardB), .ZN(n69) );
  NOR2_X2 U137 ( .A1(ALUsrc_EX), .A2(forwardB), .ZN(n68) );
  INV_X1 U138 ( .A(ALUsrc_EX), .ZN(n153) );
endmodule

