// =============================================================================
// Filename: RISC_V_tb.v
// -----------------------------------------------------------------------------
// This file exports the testbench for RISC_V.
// =============================================================================

`timescale 1 ns / 1 ps

module RISC_V_tb;
localparam CLK_PERIOD = 200;  // clock period: 200ns
// ----------------------------------
// Interface of the module
// ----------------------------------
reg		[31:0]	in;
reg 			clk;
wire    [31:0] outputdata;


// ----------------------------------
// Instantiate the module
// ----------------------------------
RISC_V uut (
	.in(in),
	.clk(clk),
	.alu_output_data(outputdata)
);


// ----------------------------------
// Clock generation
// ------------------------./----------
initial begin
  clk = 1'b0;
  forever #(CLK_PERIOD/2.0) clk = ~clk;
end



// ----------------------------------
// Input stimulus
// ----------------------------------
initial begin



in = 32'b0000_00000000_00000_000_00000_0010000;  #(CLK_PERIOD); 


in = 32'b0000_00000001_00000_000_00001_0010011;  #(CLK_PERIOD); 
in = 32'b0000_00000010_00000_000_00010_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00000011_00000_000_00011_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00000100_00000_000_00100_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00000101_00000_000_00101_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00000110_00000_000_00110_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00000111_00000_000_00111_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00001000_00000_000_01000_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00001001_00000_000_01001_0010011;  #(CLK_PERIOD); 
in = 32'b0000_00001010_00000_000_01010_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00001011_00000_000_01011_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00001100_00000_000_01100_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00001101_00000_000_01101_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00001110_00000_000_01110_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00001111_00000_000_01111_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00010000_00000_000_10000_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00010001_00000_000_10001_0010011;  #(CLK_PERIOD); 
in = 32'b0000_00010010_00000_000_10010_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00010011_00000_000_10011_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00010100_00000_000_10100_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00010101_00000_000_10101_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00010110_00000_000_10110_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00010111_00000_000_10111_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00011000_00000_000_11000_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00011001_00000_000_11001_0010011;  #(CLK_PERIOD); 
in = 32'b0000_00011010_00000_000_11010_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00011011_00000_000_11011_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00011100_00000_000_11100_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00011101_00000_000_11101_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00011110_00000_000_11110_0010011;	 #(CLK_PERIOD); 
in = 32'b0000_00011111_00000_000_11111_0010011;	 #(CLK_PERIOD);   



/*
in = 32'b0000000_00101_00000_000_00001_0010011;  #(CLK_PERIOD); 
in = 32'b0000000_00110_00000_000_00010_0010011;  #(CLK_PERIOD); 
in = 32'b0000000_00010_00001_000_00011_0110011;  #(CLK_PERIOD); 
in = 32'b0100000_00010_00011_000_00100_0110011;  #(CLK_PERIOD); 
in = 32'b0000001_00000_00010_100_00101_0010011;  #(CLK_PERIOD); 
in = 32'b0011101_10111_00001_110_00110_0010011;  #(CLK_PERIOD); 
in = 32'b0011100_11011_00110_111_00111_0010011;  #(CLK_PERIOD); 
in = 32'b0000000_00110_00101_110_01000_0110011;  #(CLK_PERIOD); 
in = 32'b0000000_00111_00110_111_01001_0110011;  #(CLK_PERIOD); 
in = 32'b0000000_00111_00101_100_01010_0110011;  #(CLK_PERIOD); 
in = 32'b0000000_00010_00001_001_01011_0110011;  #(CLK_PERIOD); 
in = 32'b0000000_00001_00010_001_01100_0010011;  #(CLK_PERIOD); 
in = 32'b0100000_00001_00110_101_01101_0110011;  #(CLK_PERIOD); 
in = 32'b0100000_00001_00110_101_01110_0010011;  #(CLK_PERIOD); 
in = 32'b0000000_00010_00001_010_01111_0110011;  #(CLK_PERIOD); 
in = 32'b0000000_00101_00001_011_10000_0010011;  #(CLK_PERIOD); 
in = 32'b0100000_01111_00010_000_00010_0110011;  #(CLK_PERIOD); 
in = 32'b1111111_00100_00010_000_11101_1100011;  #(CLK_PERIOD); 
in = 32'b0000000_00100_00010_001_00100_1100011;  #(CLK_PERIOD); 
in = 32'b0000000_00000_00001_100_10001_0110111;  #(CLK_PERIOD); 
in = 32'b0000000_00000_00000_100_00000_0010111;  #(CLK_PERIOD); 
in = 32'b0000000_11100_00000_000_10010_0010011;  #(CLK_PERIOD); 
in = 32'b0000000_11101_00000_000_10010_0010011;  #(CLK_PERIOD); 


*/










	//--------------------------------------------R_type-------------------------------------------------------------------------------------------------------

in = 32'b0000000_01100_10100_000_00101_0110011;	//1 add x5, x20,x12		x5 = 32
#(CLK_PERIOD); 

in = 32'b0100000_01100_10100_000_00110_0110011;	//2 sub x6, x20,x12		x6 = 8
#(CLK_PERIOD); 

in = 32'b0000000_01100_10100_111_00111_0110011;	//3 and x7, x20,x12     x7 = 4   0000_00010100 &  =>0000_00000100 
#(CLK_PERIOD); 									//							  	 0000_00001100

in = 32'b0000000_01100_10100_110_01000_0110011;	//4 or  x8, x20,x12     x8 = 28  0000_00010100 or =>0000_00011100
#(CLK_PERIOD);                                  //                               0000_00001100

in = 32'b0000000_01100_10100_100_01001_0110011;	//5 xor x9, x20,x12     x9 =24   0000_00010100 xor=>0000_00011000
#(CLK_PERIOD);									//                               0000_00001100

in = 32'b0000000_00100_10100_001_01010_0110011;	//6 sll x10,x20,x4      x10 =320	0000_0001_0100 <-4 0001_0100_0000
#(CLK_PERIOD); 

in = 32'b0000000_00100_10100_010_01011_0110011;	//7 slt x11,x20,x4      x11 =0	 20>4 
#(CLK_PERIOD); 

in = 32'b0100000_10100_00100_011_01100_0110011;	//8 sltu x12,x4,x20     x12= 1   4<20
#(CLK_PERIOD);

in = 32'b0000000_01100_10100_000_00000_0110011;	//9 add x0, x20,x12 	x0 = 0  register0 cannot be written
#(CLK_PERIOD); 
		
	//--------------------------------------------I_type_Imm-----------------------------------------------------------------------------------------------	

in = 32'b0000_00010000_10100_000_00000_0010011;	//10 addi x0,x20,16     x0 = 0	register0 cannot be written
#(CLK_PERIOD); 

in = 32'b0000_00010000_10100_000_00101_0010011;	//11 addi x5,x20,16		x5 = 36 
#(CLK_PERIOD); 

in = 32'b0000_00010000_10100_111_00110_0010011;	//12 andi x6,x20,16		x6 = 16   0000_00010100 & = 0000_00010000
#(CLK_PERIOD); 									//								  0000_00010000

in = 32'b0000_00010000_10100_110_00111_0010011;	//13 ori  x7,x20,16		x7 = 20	  0000_00010100 or = 0000_00010100
#(CLK_PERIOD);                                  //                                0000_00010000
 
in = 32'b0000_00010000_10100_100_01000_0010011;	//14 xori x8,x20,16		x8 = 4	  0000_00010100 xor = 0000_00000100
#(CLK_PERIOD);                                  //                                0000_00010000

in = 32'b0000000_01000_10100_001_01001_0010011;	//15 slli x9,x20,8		x9 = 5120 0000_0000_0001_0100 <- 8 0001_0100_0000_0000
#(CLK_PERIOD); 

in = 32'b1111111_11000_10100_010_01010_0010011;	//16 slti x10,x20,-8	x10 = 0  20>-8 
#(CLK_PERIOD); 

in = 32'b1111111_11000_10100_011_01011_0010011;	//17 sltiu x11,x20,-8	x11 = 1  20<unsigned(-8)
#(CLK_PERIOD); 


		
//------------------------------------------------test for data hazard	-------------------------------------------------------------------------------------------------

in = 32'b0000_00000101_00000_000_00101_0010011;	//18 addi x5,x0,5		x5 = 5  
#(CLK_PERIOD); 

in = 32'b0000000_00001_00101_000_00110_0110011;	//19 add  x6,x5,x1		x6 = 6  data hazard error:(x5 = 36, x6 = 36+1 = 37) 
#(CLK_PERIOD);                                                                  
                                                                                
in = 32'b0000_00000001_00110_000_00111_0010011;	//20 addi x7,x6,1		x7 = 7	data hazard error:(x6 =16, x7= 16+1 =17)
#(CLK_PERIOD);                                                                  
                                                                                
in = 32'b0100000_00111_01111_000_01000_0110011;	//21 sub  x8,x15,x7		x8 = 8	data hazard error :(x7 =20, x8 =15 -20 =-5)
#(CLK_PERIOD); 
		
//TEST FOR A/L RIGHT SHIFT	-------------------------------------------------------------------------

in = 32'b1111_10011100_00000_000_01010_0010011;	//22 addi x10,x0,-100   x10 = -100   (1111_10011100)
#(CLK_PERIOD); 	

//i-type
in = 32'b0000000_01000_01010_101_01011_0010011;	//23 srli x11,x10,8     x11 = 16777215 (00FF_FFFF) 	
#(CLK_PERIOD); 	      //  (-100) 1111_1111_1001_1100 ->8(Logic) =>  0000_0000_1111_1111_1111_1111_1111_1111 =00FF_FFFF


in = 32'b0100000_01000_01010_101_01100_0010011;	//24 srai x12,x10,8     x12 = -1 			
#(CLK_PERIOD); 	                            //  (-100) 1111_1111_10011100 ->8(arithmetic) =>1111_1111_1111_1111_1111_1111_1111_1111	                     								
												

//R-type
in = 32'b0000000_00100_01010_101_01101_0110011;	//25 srl x13,x10,x4     x13 =268435449	 
#(CLK_PERIOD); 									//	(-100) 1111_1111_1111_1111_1111_1111_1001_1100 ->4(Logic) 0000_1111_1111_1111_1111_1111_1111_1001					


in = 32'b0100000_00100_01010_101_01110_0110011;	//26 sra x14,x10,x4     x14= -7  (-100) 1111_1111_1001_1100 ->4(arithmetic)1111_1111_1111_1111_1111_1111_1111_1001
#(CLK_PERIOD); 

//lui
in = 32'b1111_1111_1111_1111_1111_01111_0110111;// 27 lui x15,0xFFFFF  X15 = 0XFFFFF000



 #(4*CLK_PERIOD);



$finish;
end

endmodule
